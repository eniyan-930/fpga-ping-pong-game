`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.01.2025 18:28:39
// Design Name: 
// Module Name: save_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module save_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
13'b0000000000001: color_data = 12'b111100010001;
		13'b0000000000010: color_data = 12'b111100010001;
		13'b0000000000011: color_data = 12'b111100010001;
		13'b0000000000100: color_data = 12'b111100010001;
		13'b0000000110101: color_data = 12'b111100010001;
		13'b0000001000011: color_data = 12'b111100010001;
		13'b0000001001000: color_data = 12'b111100010001;
		13'b0000001011011: color_data = 12'b111100010001;
		13'b0000001111011: color_data = 12'b111100010001;
		13'b0000010000001: color_data = 12'b111100010001;
		13'b0000010010110: color_data = 12'b111100010001;
		13'b0000100000001: color_data = 12'b111100010001;
		13'b0000100000010: color_data = 12'b111100010001;
		13'b0000100000011: color_data = 12'b111100010001;
		13'b0000100000100: color_data = 12'b111100010001;
		13'b0000100110101: color_data = 12'b111100010001;
		13'b0000101000011: color_data = 12'b111100010001;
		13'b0000101001000: color_data = 12'b111100010001;
		13'b0000101011011: color_data = 12'b111100010001;
		13'b0000101111011: color_data = 12'b111100010001;
		13'b0000110000001: color_data = 12'b111100010001;
		13'b0000110010110: color_data = 12'b111100010001;
		13'b0001000000001: color_data = 12'b111100010001;
		13'b0001000000010: color_data = 12'b111100010001;
		13'b0001000000011: color_data = 12'b111100010001;
		13'b0001000000100: color_data = 12'b111100010001;
		13'b0001000110101: color_data = 12'b111100010001;
		13'b0001001000011: color_data = 12'b111100010001;
		13'b0001001001000: color_data = 12'b111100010001;
		13'b0001001011011: color_data = 12'b111100010001;
		13'b0001001111011: color_data = 12'b111100010001;
		13'b0001010000001: color_data = 12'b111100010001;
		13'b0001010010110: color_data = 12'b111100010001;
		13'b0001100000001: color_data = 12'b111100010001;
		13'b0001100000101: color_data = 12'b111100010001;
		13'b0001100110101: color_data = 12'b111100010001;
		13'b0001101000011: color_data = 12'b111100010001;
		13'b0001101001000: color_data = 12'b111100010001;
		13'b0001101011011: color_data = 12'b111100010001;
		13'b0001101111011: color_data = 12'b111100010001;
		13'b0001110010110: color_data = 12'b111100010001;
		13'b0010000000001: color_data = 12'b111100010001;
		13'b0010000000101: color_data = 12'b111100010001;
		13'b0010000110101: color_data = 12'b111100010001;
		13'b0010001000011: color_data = 12'b111100010001;
		13'b0010001001000: color_data = 12'b111100010001;
		13'b0010001011011: color_data = 12'b111100010001;
		13'b0010001111011: color_data = 12'b111100010001;
		13'b0010010010110: color_data = 12'b111100010001;
		13'b0010100000001: color_data = 12'b111100010001;
		13'b0010100000101: color_data = 12'b111100010001;
		13'b0010100110101: color_data = 12'b111100010001;
		13'b0010101000011: color_data = 12'b111100010001;
		13'b0010101001000: color_data = 12'b111100010001;
		13'b0010101011011: color_data = 12'b111100010001;
		13'b0010101111011: color_data = 12'b111100010001;
		13'b0010110010110: color_data = 12'b111100010001;
		13'b0011000000001: color_data = 12'b111100010001;
		13'b0011000000101: color_data = 12'b111100010001;
		13'b0011000000111: color_data = 12'b111100010001;
		13'b0011000001001: color_data = 12'b111100010001;
		13'b0011000001010: color_data = 12'b111100010001;
		13'b0011000001101: color_data = 12'b111100010001;
		13'b0011000001110: color_data = 12'b111100010001;
		13'b0011000001111: color_data = 12'b111100010001;
		13'b0011000010011: color_data = 12'b111100010001;
		13'b0011000010100: color_data = 12'b111100010001;
		13'b0011000010101: color_data = 12'b111100010001;
		13'b0011000010110: color_data = 12'b111100010001;
		13'b0011000011001: color_data = 12'b111100010001;
		13'b0011000011010: color_data = 12'b111100010001;
		13'b0011000011011: color_data = 12'b111100010001;
		13'b0011000011100: color_data = 12'b111100010001;
		13'b0011000011101: color_data = 12'b111100010001;
		13'b0011000100010: color_data = 12'b111100010001;
		13'b0011000100011: color_data = 12'b111100010001;
		13'b0011000100100: color_data = 12'b111100010001;
		13'b0011000100111: color_data = 12'b111100010001;
		13'b0011000101001: color_data = 12'b111100010001;
		13'b0011000101010: color_data = 12'b111100010001;
		13'b0011000101101: color_data = 12'b111100010001;
		13'b0011000110001: color_data = 12'b111100010001;
		13'b0011000110101: color_data = 12'b111100010001;
		13'b0011000110110: color_data = 12'b111100010001;
		13'b0011000110111: color_data = 12'b111100010001;
		13'b0011000111000: color_data = 12'b111100010001;
		13'b0011000111011: color_data = 12'b111100010001;
		13'b0011001000000: color_data = 12'b111100010001;
		13'b0011001000010: color_data = 12'b111100010001;
		13'b0011001000011: color_data = 12'b111100010001;
		13'b0011001000100: color_data = 12'b111100010001;
		13'b0011001000101: color_data = 12'b111100010001;
		13'b0011001000111: color_data = 12'b111100010001;
		13'b0011001001000: color_data = 12'b111100010001;
		13'b0011001001001: color_data = 12'b111100010001;
		13'b0011001001010: color_data = 12'b111100010001;
		13'b0011001001101: color_data = 12'b111100010001;
		13'b0011001001110: color_data = 12'b111100010001;
		13'b0011001001111: color_data = 12'b111100010001;
		13'b0011001010010: color_data = 12'b111100010001;
		13'b0011001010100: color_data = 12'b111100010001;
		13'b0011001010101: color_data = 12'b111100010001;
		13'b0011001011010: color_data = 12'b111100010001;
		13'b0011001011011: color_data = 12'b111100010001;
		13'b0011001011100: color_data = 12'b111100010001;
		13'b0011001011101: color_data = 12'b111100010001;
		13'b0011001011110: color_data = 12'b111100010001;
		13'b0011001100001: color_data = 12'b111100010001;
		13'b0011001100010: color_data = 12'b111100010001;
		13'b0011001100011: color_data = 12'b111100010001;
		13'b0011001101010: color_data = 12'b111100010001;
		13'b0011001101011: color_data = 12'b111100010001;
		13'b0011001101100: color_data = 12'b111100010001;
		13'b0011001101111: color_data = 12'b111100010001;
		13'b0011001110000: color_data = 12'b111100010001;
		13'b0011001110001: color_data = 12'b111100010001;
		13'b0011001110100: color_data = 12'b111100010001;
		13'b0011001110110: color_data = 12'b111100010001;
		13'b0011001110111: color_data = 12'b111100010001;
		13'b0011001111010: color_data = 12'b111100010001;
		13'b0011001111011: color_data = 12'b111100010001;
		13'b0011001111100: color_data = 12'b111100010001;
		13'b0011001111101: color_data = 12'b111100010001;
		13'b0011010000000: color_data = 12'b111100010001;
		13'b0011010000001: color_data = 12'b111100010001;
		13'b0011010000011: color_data = 12'b111100010001;
		13'b0011010000101: color_data = 12'b111100010001;
		13'b0011010000110: color_data = 12'b111100010001;
		13'b0011010001001: color_data = 12'b111100010001;
		13'b0011010001101: color_data = 12'b111100010001;
		13'b0011010010000: color_data = 12'b111100010001;
		13'b0011010010001: color_data = 12'b111100010001;
		13'b0011010010010: color_data = 12'b111100010001;
		13'b0011010010110: color_data = 12'b111100010001;
		13'b0011100000001: color_data = 12'b111100010001;
		13'b0011100000101: color_data = 12'b111100010001;
		13'b0011100000111: color_data = 12'b111100010001;
		13'b0011100001001: color_data = 12'b111100010001;
		13'b0011100001010: color_data = 12'b111100010001;
		13'b0011100001101: color_data = 12'b111100010001;
		13'b0011100001110: color_data = 12'b111100010001;
		13'b0011100001111: color_data = 12'b111100010001;
		13'b0011100010011: color_data = 12'b111100010001;
		13'b0011100010100: color_data = 12'b111100010001;
		13'b0011100010101: color_data = 12'b111100010001;
		13'b0011100010110: color_data = 12'b111100010001;
		13'b0011100011001: color_data = 12'b111100010001;
		13'b0011100011010: color_data = 12'b111100010001;
		13'b0011100011011: color_data = 12'b111100010001;
		13'b0011100011100: color_data = 12'b111100010001;
		13'b0011100011101: color_data = 12'b111100010001;
		13'b0011100100010: color_data = 12'b111100010001;
		13'b0011100100011: color_data = 12'b111100010001;
		13'b0011100100100: color_data = 12'b111100010001;
		13'b0011100100111: color_data = 12'b111100010001;
		13'b0011100101001: color_data = 12'b111100010001;
		13'b0011100101010: color_data = 12'b111100010001;
		13'b0011100101101: color_data = 12'b111100010001;
		13'b0011100110001: color_data = 12'b111100010001;
		13'b0011100110101: color_data = 12'b111100010001;
		13'b0011100110110: color_data = 12'b111100010001;
		13'b0011100110111: color_data = 12'b111100010001;
		13'b0011100111000: color_data = 12'b111100010001;
		13'b0011100111011: color_data = 12'b111100010001;
		13'b0011101000000: color_data = 12'b111100010001;
		13'b0011101000010: color_data = 12'b111100010001;
		13'b0011101000011: color_data = 12'b111100010001;
		13'b0011101000100: color_data = 12'b111100010001;
		13'b0011101000101: color_data = 12'b111100010001;
		13'b0011101000111: color_data = 12'b111100010001;
		13'b0011101001000: color_data = 12'b111100010001;
		13'b0011101001001: color_data = 12'b111100010001;
		13'b0011101001010: color_data = 12'b111100010001;
		13'b0011101001101: color_data = 12'b111100010001;
		13'b0011101001110: color_data = 12'b111100010001;
		13'b0011101001111: color_data = 12'b111100010001;
		13'b0011101010010: color_data = 12'b111100010001;
		13'b0011101010100: color_data = 12'b111100010001;
		13'b0011101010101: color_data = 12'b111100010001;
		13'b0011101011010: color_data = 12'b111100010001;
		13'b0011101011011: color_data = 12'b111100010001;
		13'b0011101011100: color_data = 12'b111100010001;
		13'b0011101011101: color_data = 12'b111100010001;
		13'b0011101011110: color_data = 12'b111100010001;
		13'b0011101100001: color_data = 12'b111100010001;
		13'b0011101100010: color_data = 12'b111100010001;
		13'b0011101100011: color_data = 12'b111100010001;
		13'b0011101101010: color_data = 12'b111100010001;
		13'b0011101101011: color_data = 12'b111100010001;
		13'b0011101101100: color_data = 12'b111100010001;
		13'b0011101101111: color_data = 12'b111100010001;
		13'b0011101110000: color_data = 12'b111100010001;
		13'b0011101110001: color_data = 12'b111100010001;
		13'b0011101110100: color_data = 12'b111100010001;
		13'b0011101110110: color_data = 12'b111100010001;
		13'b0011101110111: color_data = 12'b111100010001;
		13'b0011101111010: color_data = 12'b111100010001;
		13'b0011101111011: color_data = 12'b111100010001;
		13'b0011101111100: color_data = 12'b111100010001;
		13'b0011101111101: color_data = 12'b111100010001;
		13'b0011110000000: color_data = 12'b111100010001;
		13'b0011110000001: color_data = 12'b111100010001;
		13'b0011110000011: color_data = 12'b111100010001;
		13'b0011110000101: color_data = 12'b111100010001;
		13'b0011110000110: color_data = 12'b111100010001;
		13'b0011110001001: color_data = 12'b111100010001;
		13'b0011110001101: color_data = 12'b111100010001;
		13'b0011110010000: color_data = 12'b111100010001;
		13'b0011110010001: color_data = 12'b111100010001;
		13'b0011110010010: color_data = 12'b111100010001;
		13'b0011110010110: color_data = 12'b111100010001;
		13'b0100000000001: color_data = 12'b111100010001;
		13'b0100000000101: color_data = 12'b111100010001;
		13'b0100000000111: color_data = 12'b111100010001;
		13'b0100000001001: color_data = 12'b111100010001;
		13'b0100000001010: color_data = 12'b111100010001;
		13'b0100000001101: color_data = 12'b111100010001;
		13'b0100000001110: color_data = 12'b111100010001;
		13'b0100000001111: color_data = 12'b111100010001;
		13'b0100000010011: color_data = 12'b111100010001;
		13'b0100000010100: color_data = 12'b111100010001;
		13'b0100000010101: color_data = 12'b111100010001;
		13'b0100000010110: color_data = 12'b111100010001;
		13'b0100000011001: color_data = 12'b111100010001;
		13'b0100000011010: color_data = 12'b111100010001;
		13'b0100000011011: color_data = 12'b111100010001;
		13'b0100000011100: color_data = 12'b111100010001;
		13'b0100000011101: color_data = 12'b111100010001;
		13'b0100000100010: color_data = 12'b111100010001;
		13'b0100000100011: color_data = 12'b111100010001;
		13'b0100000100100: color_data = 12'b111100010001;
		13'b0100000100111: color_data = 12'b111100010001;
		13'b0100000101001: color_data = 12'b111100010001;
		13'b0100000101010: color_data = 12'b111100010001;
		13'b0100000101101: color_data = 12'b111100010001;
		13'b0100000110001: color_data = 12'b111100010001;
		13'b0100000110101: color_data = 12'b111100010001;
		13'b0100000110110: color_data = 12'b111100010001;
		13'b0100000110111: color_data = 12'b111100010001;
		13'b0100000111000: color_data = 12'b111100010001;
		13'b0100000111011: color_data = 12'b111100010001;
		13'b0100001000000: color_data = 12'b111100010001;
		13'b0100001000010: color_data = 12'b111100010001;
		13'b0100001000011: color_data = 12'b111100010001;
		13'b0100001000100: color_data = 12'b111100010001;
		13'b0100001000101: color_data = 12'b111100010001;
		13'b0100001000111: color_data = 12'b111100010001;
		13'b0100001001000: color_data = 12'b111100010001;
		13'b0100001001001: color_data = 12'b111100010001;
		13'b0100001001010: color_data = 12'b111100010001;
		13'b0100001001101: color_data = 12'b111100010001;
		13'b0100001001110: color_data = 12'b111100010001;
		13'b0100001001111: color_data = 12'b111100010001;
		13'b0100001010010: color_data = 12'b111100010001;
		13'b0100001010100: color_data = 12'b111100010001;
		13'b0100001010101: color_data = 12'b111100010001;
		13'b0100001011010: color_data = 12'b111100010001;
		13'b0100001011011: color_data = 12'b111100010001;
		13'b0100001011100: color_data = 12'b111100010001;
		13'b0100001011101: color_data = 12'b111100010001;
		13'b0100001011110: color_data = 12'b111100010001;
		13'b0100001100001: color_data = 12'b111100010001;
		13'b0100001100010: color_data = 12'b111100010001;
		13'b0100001100011: color_data = 12'b111100010001;
		13'b0100001101010: color_data = 12'b111100010001;
		13'b0100001101011: color_data = 12'b111100010001;
		13'b0100001101100: color_data = 12'b111100010001;
		13'b0100001101111: color_data = 12'b111100010001;
		13'b0100001110000: color_data = 12'b111100010001;
		13'b0100001110001: color_data = 12'b111100010001;
		13'b0100001110100: color_data = 12'b111100010001;
		13'b0100001110110: color_data = 12'b111100010001;
		13'b0100001110111: color_data = 12'b111100010001;
		13'b0100001111010: color_data = 12'b111100010001;
		13'b0100001111011: color_data = 12'b111100010001;
		13'b0100001111100: color_data = 12'b111100010001;
		13'b0100001111101: color_data = 12'b111100010001;
		13'b0100010000000: color_data = 12'b111100010001;
		13'b0100010000001: color_data = 12'b111100010001;
		13'b0100010000011: color_data = 12'b111100010001;
		13'b0100010000101: color_data = 12'b111100010001;
		13'b0100010000110: color_data = 12'b111100010001;
		13'b0100010001001: color_data = 12'b111100010001;
		13'b0100010001101: color_data = 12'b111100010001;
		13'b0100010010000: color_data = 12'b111100010001;
		13'b0100010010001: color_data = 12'b111100010001;
		13'b0100010010010: color_data = 12'b111100010001;
		13'b0100010010110: color_data = 12'b111100010001;
		13'b0100100000001: color_data = 12'b111100010001;
		13'b0100100000101: color_data = 12'b111100010001;
		13'b0100100000111: color_data = 12'b111100010001;
		13'b0100100001000: color_data = 12'b111100010001;
		13'b0100100001100: color_data = 12'b111100010001;
		13'b0100100010000: color_data = 12'b111100010001;
		13'b0100100010010: color_data = 12'b111100010001;
		13'b0100100011000: color_data = 12'b111100010001;
		13'b0100100100101: color_data = 12'b111100010001;
		13'b0100100100111: color_data = 12'b111100010001;
		13'b0100100101000: color_data = 12'b111100010001;
		13'b0100100101011: color_data = 12'b111100010001;
		13'b0100100101101: color_data = 12'b111100010001;
		13'b0100100101111: color_data = 12'b111100010001;
		13'b0100100110000: color_data = 12'b111100010001;
		13'b0100100110001: color_data = 12'b111100010001;
		13'b0100100110101: color_data = 12'b111100010001;
		13'b0100100111001: color_data = 12'b111100010001;
		13'b0100100111011: color_data = 12'b111100010001;
		13'b0100101000000: color_data = 12'b111100010001;
		13'b0100101000011: color_data = 12'b111100010001;
		13'b0100101001000: color_data = 12'b111100010001;
		13'b0100101001100: color_data = 12'b111100010001;
		13'b0100101010000: color_data = 12'b111100010001;
		13'b0100101010010: color_data = 12'b111100010001;
		13'b0100101010011: color_data = 12'b111100010001;
		13'b0100101010110: color_data = 12'b111100010001;
		13'b0100101011011: color_data = 12'b111100010001;
		13'b0100101100000: color_data = 12'b111100010001;
		13'b0100101100100: color_data = 12'b111100010001;
		13'b0100101101001: color_data = 12'b111100010001;
		13'b0100101101110: color_data = 12'b111100010001;
		13'b0100101110010: color_data = 12'b111100010001;
		13'b0100101110100: color_data = 12'b111100010001;
		13'b0100101110101: color_data = 12'b111100010001;
		13'b0100101111000: color_data = 12'b111100010001;
		13'b0100101111011: color_data = 12'b111100010001;
		13'b0100110000001: color_data = 12'b111100010001;
		13'b0100110000011: color_data = 12'b111100010001;
		13'b0100110000100: color_data = 12'b111100010001;
		13'b0100110000111: color_data = 12'b111100010001;
		13'b0100110001001: color_data = 12'b111100010001;
		13'b0100110001101: color_data = 12'b111100010001;
		13'b0100110001111: color_data = 12'b111100010001;
		13'b0100110010011: color_data = 12'b111100010001;
		13'b0100110010110: color_data = 12'b111100010001;
		13'b0101000000001: color_data = 12'b111100010001;
		13'b0101000000101: color_data = 12'b111100010001;
		13'b0101000000111: color_data = 12'b111100010001;
		13'b0101000001000: color_data = 12'b111100010001;
		13'b0101000001100: color_data = 12'b111100010001;
		13'b0101000010000: color_data = 12'b111100010001;
		13'b0101000010010: color_data = 12'b111100010001;
		13'b0101000011000: color_data = 12'b111100010001;
		13'b0101000100101: color_data = 12'b111100010001;
		13'b0101000100111: color_data = 12'b111100010001;
		13'b0101000101000: color_data = 12'b111100010001;
		13'b0101000101011: color_data = 12'b111100010001;
		13'b0101000101101: color_data = 12'b111100010001;
		13'b0101000110001: color_data = 12'b111100010001;
		13'b0101000110101: color_data = 12'b111100010001;
		13'b0101000111001: color_data = 12'b111100010001;
		13'b0101000111011: color_data = 12'b111100010001;
		13'b0101001000000: color_data = 12'b111100010001;
		13'b0101001000011: color_data = 12'b111100010001;
		13'b0101001001000: color_data = 12'b111100010001;
		13'b0101001001100: color_data = 12'b111100010001;
		13'b0101001010000: color_data = 12'b111100010001;
		13'b0101001010010: color_data = 12'b111100010001;
		13'b0101001010011: color_data = 12'b111100010001;
		13'b0101001010110: color_data = 12'b111100010001;
		13'b0101001011011: color_data = 12'b111100010001;
		13'b0101001100000: color_data = 12'b111100010001;
		13'b0101001100100: color_data = 12'b111100010001;
		13'b0101001101001: color_data = 12'b111100010001;
		13'b0101001101110: color_data = 12'b111100010001;
		13'b0101001110010: color_data = 12'b111100010001;
		13'b0101001110100: color_data = 12'b111100010001;
		13'b0101001110101: color_data = 12'b111100010001;
		13'b0101001111000: color_data = 12'b111100010001;
		13'b0101001111011: color_data = 12'b111100010001;
		13'b0101010000001: color_data = 12'b111100010001;
		13'b0101010000011: color_data = 12'b111100010001;
		13'b0101010000100: color_data = 12'b111100010001;
		13'b0101010000111: color_data = 12'b111100010001;
		13'b0101010001001: color_data = 12'b111100010001;
		13'b0101010001101: color_data = 12'b111100010001;
		13'b0101010001111: color_data = 12'b111100010001;
		13'b0101010010011: color_data = 12'b111100010001;
		13'b0101010010110: color_data = 12'b111100010001;
		13'b0101100000001: color_data = 12'b111100010001;
		13'b0101100000101: color_data = 12'b111100010001;
		13'b0101100000111: color_data = 12'b111100010001;
		13'b0101100001000: color_data = 12'b111100010001;
		13'b0101100001100: color_data = 12'b111100010001;
		13'b0101100010000: color_data = 12'b111100010001;
		13'b0101100010010: color_data = 12'b111100010001;
		13'b0101100011000: color_data = 12'b111100010001;
		13'b0101100100101: color_data = 12'b111100010001;
		13'b0101100100111: color_data = 12'b111100010001;
		13'b0101100101000: color_data = 12'b111100010001;
		13'b0101100101011: color_data = 12'b111100010001;
		13'b0101100101101: color_data = 12'b111100010001;
		13'b0101100110001: color_data = 12'b111100010001;
		13'b0101100110101: color_data = 12'b111100010001;
		13'b0101100111001: color_data = 12'b111100010001;
		13'b0101100111011: color_data = 12'b111100010001;
		13'b0101101000000: color_data = 12'b111100010001;
		13'b0101101000011: color_data = 12'b111100010001;
		13'b0101101001000: color_data = 12'b111100010001;
		13'b0101101001100: color_data = 12'b111100010001;
		13'b0101101010000: color_data = 12'b111100010001;
		13'b0101101010010: color_data = 12'b111100010001;
		13'b0101101010011: color_data = 12'b111100010001;
		13'b0101101010110: color_data = 12'b111100010001;
		13'b0101101011011: color_data = 12'b111100010001;
		13'b0101101100000: color_data = 12'b111100010001;
		13'b0101101100100: color_data = 12'b111100010001;
		13'b0101101101001: color_data = 12'b111100010001;
		13'b0101101101110: color_data = 12'b111100010001;
		13'b0101101110010: color_data = 12'b111100010001;
		13'b0101101110100: color_data = 12'b111100010001;
		13'b0101101110101: color_data = 12'b111100010001;
		13'b0101101111000: color_data = 12'b111100010001;
		13'b0101101111011: color_data = 12'b111100010001;
		13'b0101110000001: color_data = 12'b111100010001;
		13'b0101110000011: color_data = 12'b111100010001;
		13'b0101110000100: color_data = 12'b111100010001;
		13'b0101110000111: color_data = 12'b111100010001;
		13'b0101110001001: color_data = 12'b111100010001;
		13'b0101110001101: color_data = 12'b111100010001;
		13'b0101110001111: color_data = 12'b111100010001;
		13'b0101110010011: color_data = 12'b111100010001;
		13'b0101110010110: color_data = 12'b111100010001;
		13'b0110000000001: color_data = 12'b111100010001;
		13'b0110000000010: color_data = 12'b111100010001;
		13'b0110000000011: color_data = 12'b111100010001;
		13'b0110000000100: color_data = 12'b111100010001;
		13'b0110000000111: color_data = 12'b111100010001;
		13'b0110000001100: color_data = 12'b111100010001;
		13'b0110000001101: color_data = 12'b111100010001;
		13'b0110000001110: color_data = 12'b111100010001;
		13'b0110000001111: color_data = 12'b111100010001;
		13'b0110000010000: color_data = 12'b111100010001;
		13'b0110000010011: color_data = 12'b111100010001;
		13'b0110000010100: color_data = 12'b111100010001;
		13'b0110000010101: color_data = 12'b111100010001;
		13'b0110000011001: color_data = 12'b111100010001;
		13'b0110000011010: color_data = 12'b111100010001;
		13'b0110000011011: color_data = 12'b111100010001;
		13'b0110000011100: color_data = 12'b111100010001;
		13'b0110000100010: color_data = 12'b111100010001;
		13'b0110000100011: color_data = 12'b111100010001;
		13'b0110000100100: color_data = 12'b111100010001;
		13'b0110000100101: color_data = 12'b111100010001;
		13'b0110000100111: color_data = 12'b111100010001;
		13'b0110000101011: color_data = 12'b111100010001;
		13'b0110000101101: color_data = 12'b111100010001;
		13'b0110000110001: color_data = 12'b111100010001;
		13'b0110000110101: color_data = 12'b111100010001;
		13'b0110000111001: color_data = 12'b111100010001;
		13'b0110000111011: color_data = 12'b111100010001;
		13'b0110001000000: color_data = 12'b111100010001;
		13'b0110001000011: color_data = 12'b111100010001;
		13'b0110001001000: color_data = 12'b111100010001;
		13'b0110001001100: color_data = 12'b111100010001;
		13'b0110001010000: color_data = 12'b111100010001;
		13'b0110001010010: color_data = 12'b111100010001;
		13'b0110001010110: color_data = 12'b111100010001;
		13'b0110001011011: color_data = 12'b111100010001;
		13'b0110001100000: color_data = 12'b111100010001;
		13'b0110001100100: color_data = 12'b111100010001;
		13'b0110001101001: color_data = 12'b111100010001;
		13'b0110001101110: color_data = 12'b111100010001;
		13'b0110001110010: color_data = 12'b111100010001;
		13'b0110001110100: color_data = 12'b111100010001;
		13'b0110001111000: color_data = 12'b111100010001;
		13'b0110001111011: color_data = 12'b111100010001;
		13'b0110010000001: color_data = 12'b111100010001;
		13'b0110010000011: color_data = 12'b111100010001;
		13'b0110010000111: color_data = 12'b111100010001;
		13'b0110010001001: color_data = 12'b111100010001;
		13'b0110010001101: color_data = 12'b111100010001;
		13'b0110010001111: color_data = 12'b111100010001;
		13'b0110010010000: color_data = 12'b111100010001;
		13'b0110010010001: color_data = 12'b111100010001;
		13'b0110010010010: color_data = 12'b111100010001;
		13'b0110010010011: color_data = 12'b111100010001;
		13'b0110010010110: color_data = 12'b111100010001;
		13'b0110100000001: color_data = 12'b111100010001;
		13'b0110100000010: color_data = 12'b111100010001;
		13'b0110100000011: color_data = 12'b111100010001;
		13'b0110100000100: color_data = 12'b111100010001;
		13'b0110100000111: color_data = 12'b111100010001;
		13'b0110100001100: color_data = 12'b111100010001;
		13'b0110100001101: color_data = 12'b111100010001;
		13'b0110100001110: color_data = 12'b111100010001;
		13'b0110100001111: color_data = 12'b111100010001;
		13'b0110100010000: color_data = 12'b111100010001;
		13'b0110100010011: color_data = 12'b111100010001;
		13'b0110100010100: color_data = 12'b111100010001;
		13'b0110100010101: color_data = 12'b111100010001;
		13'b0110100011001: color_data = 12'b111100010001;
		13'b0110100011010: color_data = 12'b111100010001;
		13'b0110100011011: color_data = 12'b111100010001;
		13'b0110100011100: color_data = 12'b111100010001;
		13'b0110100100010: color_data = 12'b111100010001;
		13'b0110100100011: color_data = 12'b111100010001;
		13'b0110100100100: color_data = 12'b111100010001;
		13'b0110100100101: color_data = 12'b111100010001;
		13'b0110100100111: color_data = 12'b111100010001;
		13'b0110100101011: color_data = 12'b111100010001;
		13'b0110100101101: color_data = 12'b111100010001;
		13'b0110100110001: color_data = 12'b111100010001;
		13'b0110100110101: color_data = 12'b111100010001;
		13'b0110100111001: color_data = 12'b111100010001;
		13'b0110100111011: color_data = 12'b111100010001;
		13'b0110101000000: color_data = 12'b111100010001;
		13'b0110101000011: color_data = 12'b111100010001;
		13'b0110101001000: color_data = 12'b111100010001;
		13'b0110101001100: color_data = 12'b111100010001;
		13'b0110101010000: color_data = 12'b111100010001;
		13'b0110101010010: color_data = 12'b111100010001;
		13'b0110101010110: color_data = 12'b111100010001;
		13'b0110101011011: color_data = 12'b111100010001;
		13'b0110101100000: color_data = 12'b111100010001;
		13'b0110101100100: color_data = 12'b111100010001;
		13'b0110101101001: color_data = 12'b111100010001;
		13'b0110101101110: color_data = 12'b111100010001;
		13'b0110101110010: color_data = 12'b111100010001;
		13'b0110101110100: color_data = 12'b111100010001;
		13'b0110101111000: color_data = 12'b111100010001;
		13'b0110101111011: color_data = 12'b111100010001;
		13'b0110110000001: color_data = 12'b111100010001;
		13'b0110110000011: color_data = 12'b111100010001;
		13'b0110110000111: color_data = 12'b111100010001;
		13'b0110110001001: color_data = 12'b111100010001;
		13'b0110110001101: color_data = 12'b111100010001;
		13'b0110110001111: color_data = 12'b111100010001;
		13'b0110110010000: color_data = 12'b111100010001;
		13'b0110110010001: color_data = 12'b111100010001;
		13'b0110110010010: color_data = 12'b111100010001;
		13'b0110110010011: color_data = 12'b111100010001;
		13'b0110110010110: color_data = 12'b111100010001;
		13'b0111000000001: color_data = 12'b111100010001;
		13'b0111000000111: color_data = 12'b111100010001;
		13'b0111000001100: color_data = 12'b111100010001;
		13'b0111000010110: color_data = 12'b111100010001;
		13'b0111000011101: color_data = 12'b111100010001;
		13'b0111000100001: color_data = 12'b111100010001;
		13'b0111000100101: color_data = 12'b111100010001;
		13'b0111000100111: color_data = 12'b111100010001;
		13'b0111000101011: color_data = 12'b111100010001;
		13'b0111000101101: color_data = 12'b111100010001;
		13'b0111000110001: color_data = 12'b111100010001;
		13'b0111000110101: color_data = 12'b111100010001;
		13'b0111000111001: color_data = 12'b111100010001;
		13'b0111000111011: color_data = 12'b111100010001;
		13'b0111000111111: color_data = 12'b111100010001;
		13'b0111001000000: color_data = 12'b111100010001;
		13'b0111001000011: color_data = 12'b111100010001;
		13'b0111001001000: color_data = 12'b111100010001;
		13'b0111001001100: color_data = 12'b111100010001;
		13'b0111001010000: color_data = 12'b111100010001;
		13'b0111001010010: color_data = 12'b111100010001;
		13'b0111001010110: color_data = 12'b111100010001;
		13'b0111001011011: color_data = 12'b111100010001;
		13'b0111001100000: color_data = 12'b111100010001;
		13'b0111001100100: color_data = 12'b111100010001;
		13'b0111001101001: color_data = 12'b111100010001;
		13'b0111001101110: color_data = 12'b111100010001;
		13'b0111001110010: color_data = 12'b111100010001;
		13'b0111001110100: color_data = 12'b111100010001;
		13'b0111001111000: color_data = 12'b111100010001;
		13'b0111001111011: color_data = 12'b111100010001;
		13'b0111010000001: color_data = 12'b111100010001;
		13'b0111010000011: color_data = 12'b111100010001;
		13'b0111010000111: color_data = 12'b111100010001;
		13'b0111010001001: color_data = 12'b111100010001;
		13'b0111010001100: color_data = 12'b111100010001;
		13'b0111010001101: color_data = 12'b111100010001;
		13'b0111010001111: color_data = 12'b111100010001;
		13'b0111100000001: color_data = 12'b111100010001;
		13'b0111100000111: color_data = 12'b111100010001;
		13'b0111100001100: color_data = 12'b111100010001;
		13'b0111100010110: color_data = 12'b111100010001;
		13'b0111100011101: color_data = 12'b111100010001;
		13'b0111100100001: color_data = 12'b111100010001;
		13'b0111100100101: color_data = 12'b111100010001;
		13'b0111100100111: color_data = 12'b111100010001;
		13'b0111100101011: color_data = 12'b111100010001;
		13'b0111100101101: color_data = 12'b111100010001;
		13'b0111100110001: color_data = 12'b111100010001;
		13'b0111100110101: color_data = 12'b111100010001;
		13'b0111100111001: color_data = 12'b111100010001;
		13'b0111100111011: color_data = 12'b111100010001;
		13'b0111100111111: color_data = 12'b111100010001;
		13'b0111101000000: color_data = 12'b111100010001;
		13'b0111101000011: color_data = 12'b111100010001;
		13'b0111101001000: color_data = 12'b111100010001;
		13'b0111101001100: color_data = 12'b111100010001;
		13'b0111101010000: color_data = 12'b111100010001;
		13'b0111101010010: color_data = 12'b111100010001;
		13'b0111101010110: color_data = 12'b111100010001;
		13'b0111101011011: color_data = 12'b111100010001;
		13'b0111101100000: color_data = 12'b111100010001;
		13'b0111101100100: color_data = 12'b111100010001;
		13'b0111101101001: color_data = 12'b111100010001;
		13'b0111101101110: color_data = 12'b111100010001;
		13'b0111101110010: color_data = 12'b111100010001;
		13'b0111101110100: color_data = 12'b111100010001;
		13'b0111101111000: color_data = 12'b111100010001;
		13'b0111101111011: color_data = 12'b111100010001;
		13'b0111110000001: color_data = 12'b111100010001;
		13'b0111110000011: color_data = 12'b111100010001;
		13'b0111110000111: color_data = 12'b111100010001;
		13'b0111110001001: color_data = 12'b111100010001;
		13'b0111110001100: color_data = 12'b111100010001;
		13'b0111110001101: color_data = 12'b111100010001;
		13'b0111110001111: color_data = 12'b111100010001;
		13'b1000000000001: color_data = 12'b111100010001;
		13'b1000000000111: color_data = 12'b111100010001;
		13'b1000000001100: color_data = 12'b111100010001;
		13'b1000000010110: color_data = 12'b111100010001;
		13'b1000000011101: color_data = 12'b111100010001;
		13'b1000000100001: color_data = 12'b111100010001;
		13'b1000000100101: color_data = 12'b111100010001;
		13'b1000000100111: color_data = 12'b111100010001;
		13'b1000000101011: color_data = 12'b111100010001;
		13'b1000000101101: color_data = 12'b111100010001;
		13'b1000000110001: color_data = 12'b111100010001;
		13'b1000000110101: color_data = 12'b111100010001;
		13'b1000000111001: color_data = 12'b111100010001;
		13'b1000000111011: color_data = 12'b111100010001;
		13'b1000000111111: color_data = 12'b111100010001;
		13'b1000001000000: color_data = 12'b111100010001;
		13'b1000001000011: color_data = 12'b111100010001;
		13'b1000001001000: color_data = 12'b111100010001;
		13'b1000001001100: color_data = 12'b111100010001;
		13'b1000001010000: color_data = 12'b111100010001;
		13'b1000001010010: color_data = 12'b111100010001;
		13'b1000001010110: color_data = 12'b111100010001;
		13'b1000001011011: color_data = 12'b111100010001;
		13'b1000001100000: color_data = 12'b111100010001;
		13'b1000001100100: color_data = 12'b111100010001;
		13'b1000001101001: color_data = 12'b111100010001;
		13'b1000001101110: color_data = 12'b111100010001;
		13'b1000001110010: color_data = 12'b111100010001;
		13'b1000001110100: color_data = 12'b111100010001;
		13'b1000001111000: color_data = 12'b111100010001;
		13'b1000001111011: color_data = 12'b111100010001;
		13'b1000010000001: color_data = 12'b111100010001;
		13'b1000010000011: color_data = 12'b111100010001;
		13'b1000010000111: color_data = 12'b111100010001;
		13'b1000010001001: color_data = 12'b111100010001;
		13'b1000010001100: color_data = 12'b111100010001;
		13'b1000010001101: color_data = 12'b111100010001;
		13'b1000010001111: color_data = 12'b111100010001;
		13'b1000100000001: color_data = 12'b111100010001;
		13'b1000100000111: color_data = 12'b111100010001;
		13'b1000100001101: color_data = 12'b111100010001;
		13'b1000100001110: color_data = 12'b111100010001;
		13'b1000100001111: color_data = 12'b111100010001;
		13'b1000100010010: color_data = 12'b111100010001;
		13'b1000100010011: color_data = 12'b111100010001;
		13'b1000100010100: color_data = 12'b111100010001;
		13'b1000100010101: color_data = 12'b111100010001;
		13'b1000100011000: color_data = 12'b111100010001;
		13'b1000100011001: color_data = 12'b111100010001;
		13'b1000100011010: color_data = 12'b111100010001;
		13'b1000100011011: color_data = 12'b111100010001;
		13'b1000100011100: color_data = 12'b111100010001;
		13'b1000100100010: color_data = 12'b111100010001;
		13'b1000100100011: color_data = 12'b111100010001;
		13'b1000100100100: color_data = 12'b111100010001;
		13'b1000100100101: color_data = 12'b111100010001;
		13'b1000100100111: color_data = 12'b111100010001;
		13'b1000100101011: color_data = 12'b111100010001;
		13'b1000100101110: color_data = 12'b111100010001;
		13'b1000100101111: color_data = 12'b111100010001;
		13'b1000100110000: color_data = 12'b111100010001;
		13'b1000100110001: color_data = 12'b111100010001;
		13'b1000100110101: color_data = 12'b111100010001;
		13'b1000100110110: color_data = 12'b111100010001;
		13'b1000100110111: color_data = 12'b111100010001;
		13'b1000100111000: color_data = 12'b111100010001;
		13'b1000100111100: color_data = 12'b111100010001;
		13'b1000100111101: color_data = 12'b111100010001;
		13'b1000100111110: color_data = 12'b111100010001;
		13'b1000101000000: color_data = 12'b111100010001;
		13'b1000101000100: color_data = 12'b111100010001;
		13'b1000101000101: color_data = 12'b111100010001;
		13'b1000101001001: color_data = 12'b111100010001;
		13'b1000101001010: color_data = 12'b111100010001;
		13'b1000101001101: color_data = 12'b111100010001;
		13'b1000101001110: color_data = 12'b111100010001;
		13'b1000101001111: color_data = 12'b111100010001;
		13'b1000101010010: color_data = 12'b111100010001;
		13'b1000101010110: color_data = 12'b111100010001;
		13'b1000101011100: color_data = 12'b111100010001;
		13'b1000101011101: color_data = 12'b111100010001;
		13'b1000101011110: color_data = 12'b111100010001;
		13'b1000101100001: color_data = 12'b111100010001;
		13'b1000101100010: color_data = 12'b111100010001;
		13'b1000101100011: color_data = 12'b111100010001;
		13'b1000101101010: color_data = 12'b111100010001;
		13'b1000101101011: color_data = 12'b111100010001;
		13'b1000101101100: color_data = 12'b111100010001;
		13'b1000101101111: color_data = 12'b111100010001;
		13'b1000101110000: color_data = 12'b111100010001;
		13'b1000101110001: color_data = 12'b111100010001;
		13'b1000101110100: color_data = 12'b111100010001;
		13'b1000101111000: color_data = 12'b111100010001;
		13'b1000101111100: color_data = 12'b111100010001;
		13'b1000101111101: color_data = 12'b111100010001;
		13'b1000110000001: color_data = 12'b111100010001;
		13'b1000110000011: color_data = 12'b111100010001;
		13'b1000110000111: color_data = 12'b111100010001;
		13'b1000110001010: color_data = 12'b111100010001;
		13'b1000110001011: color_data = 12'b111100010001;
		13'b1000110001101: color_data = 12'b111100010001;
		13'b1000110010000: color_data = 12'b111100010001;
		13'b1000110010001: color_data = 12'b111100010001;
		13'b1000110010010: color_data = 12'b111100010001;
		13'b1000110010110: color_data = 12'b111100010001;
		13'b1001000000001: color_data = 12'b111100010001;
		13'b1001000000111: color_data = 12'b111100010001;
		13'b1001000001101: color_data = 12'b111100010001;
		13'b1001000001110: color_data = 12'b111100010001;
		13'b1001000001111: color_data = 12'b111100010001;
		13'b1001000010010: color_data = 12'b111100010001;
		13'b1001000010011: color_data = 12'b111100010001;
		13'b1001000010100: color_data = 12'b111100010001;
		13'b1001000010101: color_data = 12'b111100010001;
		13'b1001000011000: color_data = 12'b111100010001;
		13'b1001000011001: color_data = 12'b111100010001;
		13'b1001000011010: color_data = 12'b111100010001;
		13'b1001000011011: color_data = 12'b111100010001;
		13'b1001000011100: color_data = 12'b111100010001;
		13'b1001000100010: color_data = 12'b111100010001;
		13'b1001000100011: color_data = 12'b111100010001;
		13'b1001000100100: color_data = 12'b111100010001;
		13'b1001000100101: color_data = 12'b111100010001;
		13'b1001000100111: color_data = 12'b111100010001;
		13'b1001000101011: color_data = 12'b111100010001;
		13'b1001000101110: color_data = 12'b111100010001;
		13'b1001000101111: color_data = 12'b111100010001;
		13'b1001000110000: color_data = 12'b111100010001;
		13'b1001000110001: color_data = 12'b111100010001;
		13'b1001000110101: color_data = 12'b111100010001;
		13'b1001000110110: color_data = 12'b111100010001;
		13'b1001000110111: color_data = 12'b111100010001;
		13'b1001000111000: color_data = 12'b111100010001;
		13'b1001000111100: color_data = 12'b111100010001;
		13'b1001000111101: color_data = 12'b111100010001;
		13'b1001000111110: color_data = 12'b111100010001;
		13'b1001001000000: color_data = 12'b111100010001;
		13'b1001001000100: color_data = 12'b111100010001;
		13'b1001001000101: color_data = 12'b111100010001;
		13'b1001001001001: color_data = 12'b111100010001;
		13'b1001001001010: color_data = 12'b111100010001;
		13'b1001001001101: color_data = 12'b111100010001;
		13'b1001001001110: color_data = 12'b111100010001;
		13'b1001001001111: color_data = 12'b111100010001;
		13'b1001001010010: color_data = 12'b111100010001;
		13'b1001001010110: color_data = 12'b111100010001;
		13'b1001001011100: color_data = 12'b111100010001;
		13'b1001001011101: color_data = 12'b111100010001;
		13'b1001001011110: color_data = 12'b111100010001;
		13'b1001001100001: color_data = 12'b111100010001;
		13'b1001001100010: color_data = 12'b111100010001;
		13'b1001001100011: color_data = 12'b111100010001;
		13'b1001001101010: color_data = 12'b111100010001;
		13'b1001001101011: color_data = 12'b111100010001;
		13'b1001001101100: color_data = 12'b111100010001;
		13'b1001001101111: color_data = 12'b111100010001;
		13'b1001001110000: color_data = 12'b111100010001;
		13'b1001001110001: color_data = 12'b111100010001;
		13'b1001001110100: color_data = 12'b111100010001;
		13'b1001001111000: color_data = 12'b111100010001;
		13'b1001001111100: color_data = 12'b111100010001;
		13'b1001001111101: color_data = 12'b111100010001;
		13'b1001010000001: color_data = 12'b111100010001;
		13'b1001010000011: color_data = 12'b111100010001;
		13'b1001010000111: color_data = 12'b111100010001;
		13'b1001010001010: color_data = 12'b111100010001;
		13'b1001010001011: color_data = 12'b111100010001;
		13'b1001010001101: color_data = 12'b111100010001;
		13'b1001010010000: color_data = 12'b111100010001;
		13'b1001010010001: color_data = 12'b111100010001;
		13'b1001010010010: color_data = 12'b111100010001;
		13'b1001010010110: color_data = 12'b111100010001;
		13'b1001100000001: color_data = 12'b111100010001;
		13'b1001100000111: color_data = 12'b111100010001;
		13'b1001100001101: color_data = 12'b111100010001;
		13'b1001100001110: color_data = 12'b111100010001;
		13'b1001100001111: color_data = 12'b111100010001;
		13'b1001100010010: color_data = 12'b111100010001;
		13'b1001100010011: color_data = 12'b111100010001;
		13'b1001100010100: color_data = 12'b111100010001;
		13'b1001100010101: color_data = 12'b111100010001;
		13'b1001100011000: color_data = 12'b111100010001;
		13'b1001100011001: color_data = 12'b111100010001;
		13'b1001100011010: color_data = 12'b111100010001;
		13'b1001100011011: color_data = 12'b111100010001;
		13'b1001100011100: color_data = 12'b111100010001;
		13'b1001100100010: color_data = 12'b111100010001;
		13'b1001100100011: color_data = 12'b111100010001;
		13'b1001100100100: color_data = 12'b111100010001;
		13'b1001100100101: color_data = 12'b111100010001;
		13'b1001100100111: color_data = 12'b111100010001;
		13'b1001100101011: color_data = 12'b111100010001;
		13'b1001100101110: color_data = 12'b111100010001;
		13'b1001100101111: color_data = 12'b111100010001;
		13'b1001100110000: color_data = 12'b111100010001;
		13'b1001100110001: color_data = 12'b111100010001;
		13'b1001100110101: color_data = 12'b111100010001;
		13'b1001100110110: color_data = 12'b111100010001;
		13'b1001100110111: color_data = 12'b111100010001;
		13'b1001100111000: color_data = 12'b111100010001;
		13'b1001100111100: color_data = 12'b111100010001;
		13'b1001100111101: color_data = 12'b111100010001;
		13'b1001100111110: color_data = 12'b111100010001;
		13'b1001101000000: color_data = 12'b111100010001;
		13'b1001101000100: color_data = 12'b111100010001;
		13'b1001101000101: color_data = 12'b111100010001;
		13'b1001101001001: color_data = 12'b111100010001;
		13'b1001101001010: color_data = 12'b111100010001;
		13'b1001101001101: color_data = 12'b111100010001;
		13'b1001101001110: color_data = 12'b111100010001;
		13'b1001101001111: color_data = 12'b111100010001;
		13'b1001101010010: color_data = 12'b111100010001;
		13'b1001101010110: color_data = 12'b111100010001;
		13'b1001101011100: color_data = 12'b111100010001;
		13'b1001101011101: color_data = 12'b111100010001;
		13'b1001101011110: color_data = 12'b111100010001;
		13'b1001101100001: color_data = 12'b111100010001;
		13'b1001101100010: color_data = 12'b111100010001;
		13'b1001101100011: color_data = 12'b111100010001;
		13'b1001101101010: color_data = 12'b111100010001;
		13'b1001101101011: color_data = 12'b111100010001;
		13'b1001101101100: color_data = 12'b111100010001;
		13'b1001101101111: color_data = 12'b111100010001;
		13'b1001101110000: color_data = 12'b111100010001;
		13'b1001101110001: color_data = 12'b111100010001;
		13'b1001101110100: color_data = 12'b111100010001;
		13'b1001101111000: color_data = 12'b111100010001;
		13'b1001101111100: color_data = 12'b111100010001;
		13'b1001101111101: color_data = 12'b111100010001;
		13'b1001110000001: color_data = 12'b111100010001;
		13'b1001110000011: color_data = 12'b111100010001;
		13'b1001110000111: color_data = 12'b111100010001;
		13'b1001110001010: color_data = 12'b111100010001;
		13'b1001110001011: color_data = 12'b111100010001;
		13'b1001110001101: color_data = 12'b111100010001;
		13'b1001110010000: color_data = 12'b111100010001;
		13'b1001110010001: color_data = 12'b111100010001;
		13'b1001110010010: color_data = 12'b111100010001;
		13'b1001110010110: color_data = 12'b111100010001;
		13'b1010000110001: color_data = 12'b111100010001;
		13'b1010100110001: color_data = 12'b111100010001;
		13'b1011000110001: color_data = 12'b111100010001;
		13'b1011100101110: color_data = 12'b111100010001;
		13'b1011100101111: color_data = 12'b111100010001;
		13'b1011100110000: color_data = 12'b111100010001;

		default: color_data = 12'b000000000000;
	endcase
endmodule
