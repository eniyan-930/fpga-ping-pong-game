module pong_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [8:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [8:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
    
		16'b0000000000001101: color_data = 12'b001110100111;
		16'b0000000000001110: color_data = 12'b001110100111;
		16'b0000000000001111: color_data = 12'b001110100111;
		16'b0000000000010000: color_data = 12'b001110100111;
		16'b0000000000010001: color_data = 12'b001110100111;
		16'b0000000000010010: color_data = 12'b001110100111;
		16'b0000000000010011: color_data = 12'b001110100111;
		16'b0000000000010100: color_data = 12'b001110100111;
		16'b0000000000010101: color_data = 12'b001110100111;
		16'b0000000000010110: color_data = 12'b001110100111;
		16'b0000000000010111: color_data = 12'b001110100111;
		16'b0000000000011000: color_data = 12'b001110100111;
		16'b0000000000011001: color_data = 12'b001110100111;
		16'b0000000000011010: color_data = 12'b001110100111;
		16'b0000000000011011: color_data = 12'b001110100111;
		16'b0000000000011100: color_data = 12'b001110100111;
		16'b0000000000011101: color_data = 12'b001110100111;
		16'b0000000000011110: color_data = 12'b001110100111;
		16'b0000000000011111: color_data = 12'b001110100111;
		16'b0000000000100000: color_data = 12'b001110100111;
		16'b0000000000100001: color_data = 12'b001110100111;
		16'b0000000000100010: color_data = 12'b001110100111;
		16'b0000000000100011: color_data = 12'b001110100111;
		16'b0000000000100100: color_data = 12'b001110100111;
		16'b0000000000101011: color_data = 12'b001110100111;
		16'b0000000000101100: color_data = 12'b001110100111;
		16'b0000000000101101: color_data = 12'b001110100111;
		16'b0000000000101110: color_data = 12'b001110100111;
		16'b0000000000101111: color_data = 12'b001110100111;
		16'b0000000000110000: color_data = 12'b001110100111;
		16'b0000000000110001: color_data = 12'b001110100111;
		16'b0000000000110010: color_data = 12'b001110100111;
		16'b0000000000110011: color_data = 12'b001110100111;
		16'b0000000000110100: color_data = 12'b001110100111;
		16'b0000000000110101: color_data = 12'b001110100111;
		16'b0000000000110110: color_data = 12'b001110100111;
		16'b0000000000110111: color_data = 12'b001110100111;
		16'b0000000001000100: color_data = 12'b001110100111;
		16'b0000000001000101: color_data = 12'b001110100111;
		16'b0000000001000110: color_data = 12'b001110100111;
		16'b0000000001000111: color_data = 12'b001110100111;
		16'b0000000001001000: color_data = 12'b001110100111;
		16'b0000000001001001: color_data = 12'b001110100111;
		16'b0000000001001010: color_data = 12'b001110100111;
		16'b0000000001001011: color_data = 12'b001110100111;
		16'b0000000001001100: color_data = 12'b001110100111;
		16'b0000000001001101: color_data = 12'b001110100111;
		16'b0000000001001110: color_data = 12'b001110100111;
		16'b0000000001001111: color_data = 12'b001110100111;
		16'b0000000001010110: color_data = 12'b001110100111;
		16'b0000000001010111: color_data = 12'b001110100111;
		16'b0000000001011000: color_data = 12'b001110100111;
		16'b0000000001011001: color_data = 12'b001110100111;
		16'b0000000001011010: color_data = 12'b001110100111;
		16'b0000000001011011: color_data = 12'b001110100111;
		16'b0000000001011100: color_data = 12'b001110100111;
		16'b0000000001011101: color_data = 12'b001110100111;
		16'b0000000001011110: color_data = 12'b001110100111;
		16'b0000000001011111: color_data = 12'b001110100111;
		16'b0000000001100000: color_data = 12'b001110100111;
		16'b0000000001100001: color_data = 12'b001110100111;
		16'b0000000001100010: color_data = 12'b001110100111;
		16'b0000000001100011: color_data = 12'b001110100111;
		16'b0000000001100100: color_data = 12'b001110100111;
		16'b0000000001100101: color_data = 12'b001110100111;
		16'b0000000001100110: color_data = 12'b001110100111;
		16'b0000000001100111: color_data = 12'b001110100111;
		16'b0000000001101000: color_data = 12'b001110100111;
		16'b0000000001101001: color_data = 12'b001110100111;
		16'b0000000001101010: color_data = 12'b001110100111;
		16'b0000000001101011: color_data = 12'b001110100111;
		16'b0000000001101100: color_data = 12'b001110100111;
		16'b0000000001101101: color_data = 12'b001110100111;
		16'b0000000001101110: color_data = 12'b001110100111;
		16'b0000000001110101: color_data = 12'b001110100111;
		16'b0000000001110110: color_data = 12'b001110100111;
		16'b0000000001110111: color_data = 12'b001110100111;
		16'b0000000001111000: color_data = 12'b001110100111;
		16'b0000000001111001: color_data = 12'b001110100111;
		16'b0000000001111010: color_data = 12'b001110100111;
		16'b0000000001111011: color_data = 12'b001110100111;
		16'b0000000001111100: color_data = 12'b001110100111;
		16'b0000000001111101: color_data = 12'b001110100111;
		16'b0000000001111110: color_data = 12'b001110100111;
		16'b0000000001111111: color_data = 12'b001110100111;
		16'b0000000010000000: color_data = 12'b001110100111;
		16'b0000000010000001: color_data = 12'b001110100111;
		16'b0000000010000010: color_data = 12'b001110100111;
		16'b0000000010000011: color_data = 12'b001110100111;
		16'b0000000010000100: color_data = 12'b001110100111;
		16'b0000000010000101: color_data = 12'b001110100111;
		16'b0000000010000110: color_data = 12'b001110100111;
		16'b0000000010000111: color_data = 12'b001110100111;
		16'b0000000010001000: color_data = 12'b001110100111;
		16'b0000000010001001: color_data = 12'b001110100111;
		16'b0000000010001010: color_data = 12'b001110100111;
		16'b0000000010001011: color_data = 12'b001110100111;
		16'b0000000010001100: color_data = 12'b001110100111;
		16'b0000000010101100: color_data = 12'b001110100111;
		16'b0000000010101101: color_data = 12'b001110100111;
		16'b0000000010101110: color_data = 12'b001110100111;
		16'b0000000010101111: color_data = 12'b001110100111;
		16'b0000000010110000: color_data = 12'b001110100111;
		16'b0000000010110001: color_data = 12'b001110100111;
		16'b0000000010110010: color_data = 12'b001110100111;
		16'b0000000010110011: color_data = 12'b001110100111;
		16'b0000000010110100: color_data = 12'b001110100111;
		16'b0000000010110101: color_data = 12'b001110100111;
		16'b0000000010110110: color_data = 12'b001110100111;
		16'b0000000010110111: color_data = 12'b001110100111;
		16'b0000000010111000: color_data = 12'b001110100111;
		16'b0000000010111001: color_data = 12'b001110100111;
		16'b0000000010111010: color_data = 12'b001110100111;
		16'b0000000010111011: color_data = 12'b001110100111;
		16'b0000000010111100: color_data = 12'b001110100111;
		16'b0000000010111101: color_data = 12'b001110100111;
		16'b0000000010111110: color_data = 12'b001110100111;
		16'b0000000010111111: color_data = 12'b001110100111;
		16'b0000000011000000: color_data = 12'b001110100111;
		16'b0000000011000001: color_data = 12'b001110100111;
		16'b0000000011000010: color_data = 12'b001110100111;
		16'b0000000011000011: color_data = 12'b001110100111;
		16'b0000000011000100: color_data = 12'b001110100111;
		16'b0000000011001011: color_data = 12'b001110100111;
		16'b0000000011001100: color_data = 12'b001110100111;
		16'b0000000011001101: color_data = 12'b001110100111;
		16'b0000000011001110: color_data = 12'b001110100111;
		16'b0000000011001111: color_data = 12'b001110100111;
		16'b0000000011010000: color_data = 12'b001110100111;
		16'b0000000011010001: color_data = 12'b001110100111;
		16'b0000000011010010: color_data = 12'b001110100111;
		16'b0000000011010011: color_data = 12'b001110100111;
		16'b0000000011010100: color_data = 12'b001110100111;
		16'b0000000011010101: color_data = 12'b001110100111;
		16'b0000000011010110: color_data = 12'b001110100111;
		16'b0000000011010111: color_data = 12'b001110100111;
		16'b0000000011011000: color_data = 12'b001110100111;
		16'b0000000011011001: color_data = 12'b001110100111;
		16'b0000000011011010: color_data = 12'b001110100111;
		16'b0000000011011011: color_data = 12'b001110100111;
		16'b0000000011011100: color_data = 12'b001110100111;
		16'b0000000011011101: color_data = 12'b001110100111;
		16'b0000000011011110: color_data = 12'b001110100111;
		16'b0000000011011111: color_data = 12'b001110100111;
		16'b0000000011100000: color_data = 12'b001110100111;
		16'b0000000011100001: color_data = 12'b001110100111;
		16'b0000000011100010: color_data = 12'b001110100111;
		16'b0000000011100011: color_data = 12'b001110100111;
		16'b0000000011100100: color_data = 12'b001110100111;
		16'b0000000011100101: color_data = 12'b001110100111;
		16'b0000000011100110: color_data = 12'b001110100111;
		16'b0000000011100111: color_data = 12'b001110100111;
		16'b0000000011101000: color_data = 12'b001110100111;
		16'b0000000011101001: color_data = 12'b001110100111;
		16'b0000000011101010: color_data = 12'b001110100111;
		16'b0000000011101011: color_data = 12'b001110100111;
		16'b0000000011101100: color_data = 12'b001110100111;
		16'b0000000011101101: color_data = 12'b001110100111;
		16'b0000000011101110: color_data = 12'b001110100111;
		16'b0000000011101111: color_data = 12'b001110100111;
		16'b0000000011111100: color_data = 12'b001110100111;
		16'b0000000011111101: color_data = 12'b001110100111;
		16'b0000000011111110: color_data = 12'b001110100111;
		16'b0000000011111111: color_data = 12'b001110100111;
		16'b0000000100000000: color_data = 12'b001110100111;
		16'b0000000100000001: color_data = 12'b001110100111;
		16'b0000000100000010: color_data = 12'b001110100111;
		16'b0000000100000011: color_data = 12'b001110100111;
		16'b0000000100000100: color_data = 12'b001110100111;
		16'b0000000100000101: color_data = 12'b001110100111;
		16'b0000000100000110: color_data = 12'b001110100111;
		16'b0000000100000111: color_data = 12'b001110100111;
		16'b0000000100001000: color_data = 12'b001110100111;
		16'b0000000100001001: color_data = 12'b001110100111;
		16'b0000000100001010: color_data = 12'b001110100111;
		16'b0000000100001011: color_data = 12'b001110100111;
		16'b0000000100001100: color_data = 12'b001110100111;
		16'b0000000100001101: color_data = 12'b001110100111;
		16'b0000000100001110: color_data = 12'b001110100111;
		16'b0000000100001111: color_data = 12'b001110100111;
		16'b0000000100010000: color_data = 12'b001110100111;
		16'b0000000100010001: color_data = 12'b001110100111;
		16'b0000000100010010: color_data = 12'b001110100111;
		16'b0000000100010011: color_data = 12'b001110100111;
		16'b0000000100010100: color_data = 12'b001110100111;
		16'b0000000100010101: color_data = 12'b001110100111;
		16'b0000000100010110: color_data = 12'b001110100111;
		16'b0000000100010111: color_data = 12'b001110100111;
		16'b0000000100011000: color_data = 12'b001110100111;
		16'b0000000100011001: color_data = 12'b001110100111;
		16'b0000000100011010: color_data = 12'b001110100111;
		16'b0000000100011011: color_data = 12'b001110100111;
		16'b0000000100011100: color_data = 12'b001110100111;
		16'b0000000100011101: color_data = 12'b001110100111;
		16'b0000000100011110: color_data = 12'b001110100111;
		16'b0000000100011111: color_data = 12'b001110100111;
		16'b0000000100100000: color_data = 12'b001110100111;
		16'b0000000100101101: color_data = 12'b001110100111;
		16'b0000000100101110: color_data = 12'b001110100111;
		16'b0000000100101111: color_data = 12'b001110100111;
		16'b0000000100110000: color_data = 12'b001110100111;
		16'b0000000100110001: color_data = 12'b001110100111;
		16'b0000000100110010: color_data = 12'b001110100111;
		16'b0000000100110011: color_data = 12'b001110100111;
		16'b0000000100110100: color_data = 12'b001110100111;
		16'b0000000100110101: color_data = 12'b001110100111;
		16'b0000000100110110: color_data = 12'b001110100111;
		16'b0000000100110111: color_data = 12'b001110100111;
		16'b0000000100111000: color_data = 12'b001110100111;
		16'b0000000100111001: color_data = 12'b001110100111;
		16'b0000000100111010: color_data = 12'b001110100111;
		16'b0000000100111011: color_data = 12'b001110100111;
		16'b0000000100111100: color_data = 12'b001110100111;
		16'b0000000100111101: color_data = 12'b001110100111;
		16'b0000000100111110: color_data = 12'b001110100111;
		16'b0000000100111111: color_data = 12'b001110100111;
		16'b0000000101000000: color_data = 12'b001110100111;
		16'b0000000101000001: color_data = 12'b001110100111;
		16'b0000000101000010: color_data = 12'b001110100111;
		16'b0000000101000011: color_data = 12'b001110100111;
		16'b0000000101000100: color_data = 12'b001110100111;
		16'b0000000101100100: color_data = 12'b001110100111;
		16'b0000000101100101: color_data = 12'b001110100111;
		16'b0000000101100110: color_data = 12'b001110100111;
		16'b0000000101100111: color_data = 12'b001110100111;
		16'b0000000101101000: color_data = 12'b001110100111;
		16'b0000000101101001: color_data = 12'b001110100111;
		16'b0000000101101010: color_data = 12'b001110100111;
		16'b0000000101101011: color_data = 12'b001110100111;
		16'b0000000101101100: color_data = 12'b001110100111;
		16'b0000000101101101: color_data = 12'b001110100111;
		16'b0000000101101110: color_data = 12'b001110100111;
		16'b0000000101101111: color_data = 12'b001110100111;
		16'b0000000101110000: color_data = 12'b001110100111;
		16'b0000000101110001: color_data = 12'b001110100111;
		16'b0000000101110010: color_data = 12'b001110100111;
		16'b0000000101110011: color_data = 12'b001110100111;
		16'b0000000101110100: color_data = 12'b001110100111;
		16'b0000000101110101: color_data = 12'b001110100111;
		16'b0000000101110110: color_data = 12'b001110100111;
		16'b0000000101110111: color_data = 12'b001110100111;
		16'b0000000101111000: color_data = 12'b001110100111;
		16'b0000000101111001: color_data = 12'b001110100111;
		16'b0000000101111010: color_data = 12'b001110100111;
		16'b0000000101111011: color_data = 12'b001110100111;
		16'b0000001000001101: color_data = 12'b001110100111;
		16'b0000001000001110: color_data = 12'b001110100111;
		16'b0000001000001111: color_data = 12'b001110100111;
		16'b0000001000010000: color_data = 12'b001110100111;
		16'b0000001000010001: color_data = 12'b001110100111;
		16'b0000001000010010: color_data = 12'b001110100111;
		16'b0000001000010011: color_data = 12'b001110100111;
		16'b0000001000010100: color_data = 12'b001110100111;
		16'b0000001000010101: color_data = 12'b001110100111;
		16'b0000001000010110: color_data = 12'b001110100111;
		16'b0000001000010111: color_data = 12'b001110100111;
		16'b0000001000011000: color_data = 12'b001110100111;
		16'b0000001000011001: color_data = 12'b001110100111;
		16'b0000001000011010: color_data = 12'b001110100111;
		16'b0000001000011011: color_data = 12'b001110100111;
		16'b0000001000011100: color_data = 12'b001110100111;
		16'b0000001000011101: color_data = 12'b001110100111;
		16'b0000001000011110: color_data = 12'b001110100111;
		16'b0000001000011111: color_data = 12'b001110100111;
		16'b0000001000100000: color_data = 12'b001110100111;
		16'b0000001000100001: color_data = 12'b001110100111;
		16'b0000001000100010: color_data = 12'b001110100111;
		16'b0000001000100011: color_data = 12'b001110100111;
		16'b0000001000100100: color_data = 12'b001110100111;
		16'b0000001000101011: color_data = 12'b001110100111;
		16'b0000001000101100: color_data = 12'b001110100111;
		16'b0000001000101101: color_data = 12'b001110100111;
		16'b0000001000101110: color_data = 12'b001110100111;
		16'b0000001000101111: color_data = 12'b001110100111;
		16'b0000001000110000: color_data = 12'b001110100111;
		16'b0000001000110001: color_data = 12'b001110100111;
		16'b0000001000110010: color_data = 12'b001110100111;
		16'b0000001000110011: color_data = 12'b001110100111;
		16'b0000001000110100: color_data = 12'b001110100111;
		16'b0000001000110101: color_data = 12'b001110100111;
		16'b0000001000110110: color_data = 12'b001110100111;
		16'b0000001000110111: color_data = 12'b001110100111;
		16'b0000001001000100: color_data = 12'b001110100111;
		16'b0000001001000101: color_data = 12'b001110100111;
		16'b0000001001000110: color_data = 12'b001110100111;
		16'b0000001001000111: color_data = 12'b001110100111;
		16'b0000001001001000: color_data = 12'b001110100111;
		16'b0000001001001001: color_data = 12'b001110100111;
		16'b0000001001001010: color_data = 12'b001110100111;
		16'b0000001001001011: color_data = 12'b001110100111;
		16'b0000001001001100: color_data = 12'b001110100111;
		16'b0000001001001101: color_data = 12'b001110100111;
		16'b0000001001001110: color_data = 12'b001110100111;
		16'b0000001001001111: color_data = 12'b001110100111;
		16'b0000001001010110: color_data = 12'b001110100111;
		16'b0000001001010111: color_data = 12'b001110100111;
		16'b0000001001011000: color_data = 12'b001110100111;
		16'b0000001001011001: color_data = 12'b001110100111;
		16'b0000001001011010: color_data = 12'b001110100111;
		16'b0000001001011011: color_data = 12'b001110100111;
		16'b0000001001011100: color_data = 12'b001110100111;
		16'b0000001001011101: color_data = 12'b001110100111;
		16'b0000001001011110: color_data = 12'b001110100111;
		16'b0000001001011111: color_data = 12'b001110100111;
		16'b0000001001100000: color_data = 12'b001110100111;
		16'b0000001001100001: color_data = 12'b001110100111;
		16'b0000001001100010: color_data = 12'b001110100111;
		16'b0000001001100011: color_data = 12'b001110100111;
		16'b0000001001100100: color_data = 12'b001110100111;
		16'b0000001001100101: color_data = 12'b001110100111;
		16'b0000001001100110: color_data = 12'b001110100111;
		16'b0000001001100111: color_data = 12'b001110100111;
		16'b0000001001101000: color_data = 12'b001110100111;
		16'b0000001001101001: color_data = 12'b001110100111;
		16'b0000001001101010: color_data = 12'b001110100111;
		16'b0000001001101011: color_data = 12'b001110100111;
		16'b0000001001101100: color_data = 12'b001110100111;
		16'b0000001001101101: color_data = 12'b001110100111;
		16'b0000001001101110: color_data = 12'b001110100111;
		16'b0000001001110101: color_data = 12'b001110100111;
		16'b0000001001110110: color_data = 12'b001110100111;
		16'b0000001001110111: color_data = 12'b001110100111;
		16'b0000001001111000: color_data = 12'b001110100111;
		16'b0000001001111001: color_data = 12'b001110100111;
		16'b0000001001111010: color_data = 12'b001110100111;
		16'b0000001001111011: color_data = 12'b001110100111;
		16'b0000001001111100: color_data = 12'b001110100111;
		16'b0000001001111101: color_data = 12'b001110100111;
		16'b0000001001111110: color_data = 12'b001110100111;
		16'b0000001001111111: color_data = 12'b001110100111;
		16'b0000001010000000: color_data = 12'b001110100111;
		16'b0000001010000001: color_data = 12'b001110100111;
		16'b0000001010000010: color_data = 12'b001110100111;
		16'b0000001010000011: color_data = 12'b001110100111;
		16'b0000001010000100: color_data = 12'b001110100111;
		16'b0000001010000101: color_data = 12'b001110100111;
		16'b0000001010000110: color_data = 12'b001110100111;
		16'b0000001010000111: color_data = 12'b001110100111;
		16'b0000001010001000: color_data = 12'b001110100111;
		16'b0000001010001001: color_data = 12'b001110100111;
		16'b0000001010001010: color_data = 12'b001110100111;
		16'b0000001010001011: color_data = 12'b001110100111;
		16'b0000001010001100: color_data = 12'b001110100111;
		16'b0000001010101100: color_data = 12'b001110100111;
		16'b0000001010101101: color_data = 12'b001110100111;
		16'b0000001010101110: color_data = 12'b001110100111;
		16'b0000001010101111: color_data = 12'b001110100111;
		16'b0000001010110000: color_data = 12'b001110100111;
		16'b0000001010110001: color_data = 12'b001110100111;
		16'b0000001010110010: color_data = 12'b001110100111;
		16'b0000001010110011: color_data = 12'b001110100111;
		16'b0000001010110100: color_data = 12'b001110100111;
		16'b0000001010110101: color_data = 12'b001110100111;
		16'b0000001010110110: color_data = 12'b001110100111;
		16'b0000001010110111: color_data = 12'b001110100111;
		16'b0000001010111000: color_data = 12'b001110100111;
		16'b0000001010111001: color_data = 12'b001110100111;
		16'b0000001010111010: color_data = 12'b001110100111;
		16'b0000001010111011: color_data = 12'b001110100111;
		16'b0000001010111100: color_data = 12'b001110100111;
		16'b0000001010111101: color_data = 12'b001110100111;
		16'b0000001010111110: color_data = 12'b001110100111;
		16'b0000001010111111: color_data = 12'b001110100111;
		16'b0000001011000000: color_data = 12'b001110100111;
		16'b0000001011000001: color_data = 12'b001110100111;
		16'b0000001011000010: color_data = 12'b001110100111;
		16'b0000001011000011: color_data = 12'b001110100111;
		16'b0000001011000100: color_data = 12'b001110100111;
		16'b0000001011001011: color_data = 12'b001110100111;
		16'b0000001011001100: color_data = 12'b001110100111;
		16'b0000001011001101: color_data = 12'b001110100111;
		16'b0000001011001110: color_data = 12'b001110100111;
		16'b0000001011001111: color_data = 12'b001110100111;
		16'b0000001011010000: color_data = 12'b001110100111;
		16'b0000001011010001: color_data = 12'b001110100111;
		16'b0000001011010010: color_data = 12'b001110100111;
		16'b0000001011010011: color_data = 12'b001110100111;
		16'b0000001011010100: color_data = 12'b001110100111;
		16'b0000001011010101: color_data = 12'b001110100111;
		16'b0000001011010110: color_data = 12'b001110100111;
		16'b0000001011010111: color_data = 12'b001110100111;
		16'b0000001011011000: color_data = 12'b001110100111;
		16'b0000001011011001: color_data = 12'b001110100111;
		16'b0000001011011010: color_data = 12'b001110100111;
		16'b0000001011011011: color_data = 12'b001110100111;
		16'b0000001011011100: color_data = 12'b001110100111;
		16'b0000001011011101: color_data = 12'b001110100111;
		16'b0000001011011110: color_data = 12'b001110100111;
		16'b0000001011011111: color_data = 12'b001110100111;
		16'b0000001011100000: color_data = 12'b001110100111;
		16'b0000001011100001: color_data = 12'b001110100111;
		16'b0000001011100010: color_data = 12'b001110100111;
		16'b0000001011100011: color_data = 12'b001110100111;
		16'b0000001011100100: color_data = 12'b001110100111;
		16'b0000001011100101: color_data = 12'b001110100111;
		16'b0000001011100110: color_data = 12'b001110100111;
		16'b0000001011100111: color_data = 12'b001110100111;
		16'b0000001011101000: color_data = 12'b001110100111;
		16'b0000001011101001: color_data = 12'b001110100111;
		16'b0000001011101010: color_data = 12'b001110100111;
		16'b0000001011101011: color_data = 12'b001110100111;
		16'b0000001011101100: color_data = 12'b001110100111;
		16'b0000001011101101: color_data = 12'b001110100111;
		16'b0000001011101110: color_data = 12'b001110100111;
		16'b0000001011101111: color_data = 12'b001110100111;
		16'b0000001011111100: color_data = 12'b001110100111;
		16'b0000001011111101: color_data = 12'b001110100111;
		16'b0000001011111110: color_data = 12'b001110100111;
		16'b0000001011111111: color_data = 12'b001110100111;
		16'b0000001100000000: color_data = 12'b001110100111;
		16'b0000001100000001: color_data = 12'b001110100111;
		16'b0000001100000010: color_data = 12'b001110100111;
		16'b0000001100000011: color_data = 12'b001110100111;
		16'b0000001100000100: color_data = 12'b001110100111;
		16'b0000001100000101: color_data = 12'b001110100111;
		16'b0000001100000110: color_data = 12'b001110100111;
		16'b0000001100000111: color_data = 12'b001110100111;
		16'b0000001100001000: color_data = 12'b001110100111;
		16'b0000001100001001: color_data = 12'b001110100111;
		16'b0000001100001010: color_data = 12'b001110100111;
		16'b0000001100001011: color_data = 12'b001110100111;
		16'b0000001100001100: color_data = 12'b001110100111;
		16'b0000001100001101: color_data = 12'b001110100111;
		16'b0000001100001110: color_data = 12'b001110100111;
		16'b0000001100001111: color_data = 12'b001110100111;
		16'b0000001100010000: color_data = 12'b001110100111;
		16'b0000001100010001: color_data = 12'b001110100111;
		16'b0000001100010010: color_data = 12'b001110100111;
		16'b0000001100010011: color_data = 12'b001110100111;
		16'b0000001100010100: color_data = 12'b001110100111;
		16'b0000001100010101: color_data = 12'b001110100111;
		16'b0000001100010110: color_data = 12'b001110100111;
		16'b0000001100010111: color_data = 12'b001110100111;
		16'b0000001100011000: color_data = 12'b001110100111;
		16'b0000001100011001: color_data = 12'b001110100111;
		16'b0000001100011010: color_data = 12'b001110100111;
		16'b0000001100011011: color_data = 12'b001110100111;
		16'b0000001100011100: color_data = 12'b001110100111;
		16'b0000001100011101: color_data = 12'b001110100111;
		16'b0000001100011110: color_data = 12'b001110100111;
		16'b0000001100011111: color_data = 12'b001110100111;
		16'b0000001100100000: color_data = 12'b001110100111;
		16'b0000001100101101: color_data = 12'b001110100111;
		16'b0000001100101110: color_data = 12'b001110100111;
		16'b0000001100101111: color_data = 12'b001110100111;
		16'b0000001100110000: color_data = 12'b001110100111;
		16'b0000001100110001: color_data = 12'b001110100111;
		16'b0000001100110010: color_data = 12'b001110100111;
		16'b0000001100110011: color_data = 12'b001110100111;
		16'b0000001100110100: color_data = 12'b001110100111;
		16'b0000001100110101: color_data = 12'b001110100111;
		16'b0000001100110110: color_data = 12'b001110100111;
		16'b0000001100110111: color_data = 12'b001110100111;
		16'b0000001100111000: color_data = 12'b001110100111;
		16'b0000001100111001: color_data = 12'b001110100111;
		16'b0000001100111010: color_data = 12'b001110100111;
		16'b0000001100111011: color_data = 12'b001110100111;
		16'b0000001100111100: color_data = 12'b001110100111;
		16'b0000001100111101: color_data = 12'b001110100111;
		16'b0000001100111110: color_data = 12'b001110100111;
		16'b0000001100111111: color_data = 12'b001110100111;
		16'b0000001101000000: color_data = 12'b001110100111;
		16'b0000001101000001: color_data = 12'b001110100111;
		16'b0000001101000010: color_data = 12'b001110100111;
		16'b0000001101000011: color_data = 12'b001110100111;
		16'b0000001101000100: color_data = 12'b001110100111;
		16'b0000001101100100: color_data = 12'b001110100111;
		16'b0000001101100101: color_data = 12'b001110100111;
		16'b0000001101100110: color_data = 12'b001110100111;
		16'b0000001101100111: color_data = 12'b001110100111;
		16'b0000001101101000: color_data = 12'b001110100111;
		16'b0000001101101001: color_data = 12'b001110100111;
		16'b0000001101101010: color_data = 12'b001110100111;
		16'b0000001101101011: color_data = 12'b001110100111;
		16'b0000001101101100: color_data = 12'b001110100111;
		16'b0000001101101101: color_data = 12'b001110100111;
		16'b0000001101101110: color_data = 12'b001110100111;
		16'b0000001101101111: color_data = 12'b001110100111;
		16'b0000001101110000: color_data = 12'b001110100111;
		16'b0000001101110001: color_data = 12'b001110100111;
		16'b0000001101110010: color_data = 12'b001110100111;
		16'b0000001101110011: color_data = 12'b001110100111;
		16'b0000001101110100: color_data = 12'b001110100111;
		16'b0000001101110101: color_data = 12'b001110100111;
		16'b0000001101110110: color_data = 12'b001110100111;
		16'b0000001101110111: color_data = 12'b001110100111;
		16'b0000001101111000: color_data = 12'b001110100111;
		16'b0000001101111001: color_data = 12'b001110100111;
		16'b0000001101111010: color_data = 12'b001110100111;
		16'b0000001101111011: color_data = 12'b001110100111;
		16'b0000010000001101: color_data = 12'b001110100111;
		16'b0000010000001110: color_data = 12'b001110100111;
		16'b0000010000001111: color_data = 12'b001110100111;
		16'b0000010000010000: color_data = 12'b001110100111;
		16'b0000010000010001: color_data = 12'b001110100111;
		16'b0000010000010010: color_data = 12'b001110100111;
		16'b0000010000010011: color_data = 12'b001110100111;
		16'b0000010000010100: color_data = 12'b001110100111;
		16'b0000010000010101: color_data = 12'b001110100111;
		16'b0000010000010110: color_data = 12'b001110100111;
		16'b0000010000010111: color_data = 12'b001110100111;
		16'b0000010000011000: color_data = 12'b001110100111;
		16'b0000010000011001: color_data = 12'b001110100111;
		16'b0000010000011010: color_data = 12'b001110100111;
		16'b0000010000011011: color_data = 12'b001110100111;
		16'b0000010000011100: color_data = 12'b001110100111;
		16'b0000010000011101: color_data = 12'b001110100111;
		16'b0000010000011110: color_data = 12'b001110100111;
		16'b0000010000011111: color_data = 12'b001110100111;
		16'b0000010000100000: color_data = 12'b001110100111;
		16'b0000010000100001: color_data = 12'b001110100111;
		16'b0000010000100010: color_data = 12'b001110100111;
		16'b0000010000100011: color_data = 12'b001110100111;
		16'b0000010000100100: color_data = 12'b001110100111;
		16'b0000010000101011: color_data = 12'b001110100111;
		16'b0000010000101100: color_data = 12'b001110100111;
		16'b0000010000101101: color_data = 12'b001110100111;
		16'b0000010000101110: color_data = 12'b001110100111;
		16'b0000010000101111: color_data = 12'b001110100111;
		16'b0000010000110000: color_data = 12'b001110100111;
		16'b0000010000110001: color_data = 12'b001110100111;
		16'b0000010000110010: color_data = 12'b001110100111;
		16'b0000010000110011: color_data = 12'b001110100111;
		16'b0000010000110100: color_data = 12'b001110100111;
		16'b0000010000110101: color_data = 12'b001110100111;
		16'b0000010000110110: color_data = 12'b001110100111;
		16'b0000010000110111: color_data = 12'b001110100111;
		16'b0000010001000100: color_data = 12'b001110100111;
		16'b0000010001000101: color_data = 12'b001110100111;
		16'b0000010001000110: color_data = 12'b001110100111;
		16'b0000010001000111: color_data = 12'b001110100111;
		16'b0000010001001000: color_data = 12'b001110100111;
		16'b0000010001001001: color_data = 12'b001110100111;
		16'b0000010001001010: color_data = 12'b001110100111;
		16'b0000010001001011: color_data = 12'b001110100111;
		16'b0000010001001100: color_data = 12'b001110100111;
		16'b0000010001001101: color_data = 12'b001110100111;
		16'b0000010001001110: color_data = 12'b001110100111;
		16'b0000010001001111: color_data = 12'b001110100111;
		16'b0000010001010110: color_data = 12'b001110100111;
		16'b0000010001010111: color_data = 12'b001110100111;
		16'b0000010001011000: color_data = 12'b001110100111;
		16'b0000010001011001: color_data = 12'b001110100111;
		16'b0000010001011010: color_data = 12'b001110100111;
		16'b0000010001011011: color_data = 12'b001110100111;
		16'b0000010001011100: color_data = 12'b001110100111;
		16'b0000010001011101: color_data = 12'b001110100111;
		16'b0000010001011110: color_data = 12'b001110100111;
		16'b0000010001011111: color_data = 12'b001110100111;
		16'b0000010001100000: color_data = 12'b001110100111;
		16'b0000010001100001: color_data = 12'b001110100111;
		16'b0000010001100010: color_data = 12'b001110100111;
		16'b0000010001100011: color_data = 12'b001110100111;
		16'b0000010001100100: color_data = 12'b001110100111;
		16'b0000010001100101: color_data = 12'b001110100111;
		16'b0000010001100110: color_data = 12'b001110100111;
		16'b0000010001100111: color_data = 12'b001110100111;
		16'b0000010001101000: color_data = 12'b001110100111;
		16'b0000010001101001: color_data = 12'b001110100111;
		16'b0000010001101010: color_data = 12'b001110100111;
		16'b0000010001101011: color_data = 12'b001110100111;
		16'b0000010001101100: color_data = 12'b001110100111;
		16'b0000010001101101: color_data = 12'b001110100111;
		16'b0000010001101110: color_data = 12'b001110100111;
		16'b0000010001110101: color_data = 12'b001110100111;
		16'b0000010001110110: color_data = 12'b001110100111;
		16'b0000010001110111: color_data = 12'b001110100111;
		16'b0000010001111000: color_data = 12'b001110100111;
		16'b0000010001111001: color_data = 12'b001110100111;
		16'b0000010001111010: color_data = 12'b001110100111;
		16'b0000010001111011: color_data = 12'b001110100111;
		16'b0000010001111100: color_data = 12'b001110100111;
		16'b0000010001111101: color_data = 12'b001110100111;
		16'b0000010001111110: color_data = 12'b001110100111;
		16'b0000010001111111: color_data = 12'b001110100111;
		16'b0000010010000000: color_data = 12'b001110100111;
		16'b0000010010000001: color_data = 12'b001110100111;
		16'b0000010010000010: color_data = 12'b001110100111;
		16'b0000010010000011: color_data = 12'b001110100111;
		16'b0000010010000100: color_data = 12'b001110100111;
		16'b0000010010000101: color_data = 12'b001110100111;
		16'b0000010010000110: color_data = 12'b001110100111;
		16'b0000010010000111: color_data = 12'b001110100111;
		16'b0000010010001000: color_data = 12'b001110100111;
		16'b0000010010001001: color_data = 12'b001110100111;
		16'b0000010010001010: color_data = 12'b001110100111;
		16'b0000010010001011: color_data = 12'b001110100111;
		16'b0000010010001100: color_data = 12'b001110100111;
		16'b0000010010101100: color_data = 12'b001110100111;
		16'b0000010010101101: color_data = 12'b001110100111;
		16'b0000010010101110: color_data = 12'b001110100111;
		16'b0000010010101111: color_data = 12'b001110100111;
		16'b0000010010110000: color_data = 12'b001110100111;
		16'b0000010010110001: color_data = 12'b001110100111;
		16'b0000010010110010: color_data = 12'b001110100111;
		16'b0000010010110011: color_data = 12'b001110100111;
		16'b0000010010110100: color_data = 12'b001110100111;
		16'b0000010010110101: color_data = 12'b001110100111;
		16'b0000010010110110: color_data = 12'b001110100111;
		16'b0000010010110111: color_data = 12'b001110100111;
		16'b0000010010111000: color_data = 12'b001110100111;
		16'b0000010010111001: color_data = 12'b001110100111;
		16'b0000010010111010: color_data = 12'b001110100111;
		16'b0000010010111011: color_data = 12'b001110100111;
		16'b0000010010111100: color_data = 12'b001110100111;
		16'b0000010010111101: color_data = 12'b001110100111;
		16'b0000010010111110: color_data = 12'b001110100111;
		16'b0000010010111111: color_data = 12'b001110100111;
		16'b0000010011000000: color_data = 12'b001110100111;
		16'b0000010011000001: color_data = 12'b001110100111;
		16'b0000010011000010: color_data = 12'b001110100111;
		16'b0000010011000011: color_data = 12'b001110100111;
		16'b0000010011000100: color_data = 12'b001110100111;
		16'b0000010011001011: color_data = 12'b001110100111;
		16'b0000010011001100: color_data = 12'b001110100111;
		16'b0000010011001101: color_data = 12'b001110100111;
		16'b0000010011001110: color_data = 12'b001110100111;
		16'b0000010011001111: color_data = 12'b001110100111;
		16'b0000010011010000: color_data = 12'b001110100111;
		16'b0000010011010001: color_data = 12'b001110100111;
		16'b0000010011010010: color_data = 12'b001110100111;
		16'b0000010011010011: color_data = 12'b001110100111;
		16'b0000010011010100: color_data = 12'b001110100111;
		16'b0000010011010101: color_data = 12'b001110100111;
		16'b0000010011010110: color_data = 12'b001110100111;
		16'b0000010011010111: color_data = 12'b001110100111;
		16'b0000010011011000: color_data = 12'b001110100111;
		16'b0000010011011001: color_data = 12'b001110100111;
		16'b0000010011011010: color_data = 12'b001110100111;
		16'b0000010011011011: color_data = 12'b001110100111;
		16'b0000010011011100: color_data = 12'b001110100111;
		16'b0000010011011101: color_data = 12'b001110100111;
		16'b0000010011011110: color_data = 12'b001110100111;
		16'b0000010011011111: color_data = 12'b001110100111;
		16'b0000010011100000: color_data = 12'b001110100111;
		16'b0000010011100001: color_data = 12'b001110100111;
		16'b0000010011100010: color_data = 12'b001110100111;
		16'b0000010011100011: color_data = 12'b001110100111;
		16'b0000010011100100: color_data = 12'b001110100111;
		16'b0000010011100101: color_data = 12'b001110100111;
		16'b0000010011100110: color_data = 12'b001110100111;
		16'b0000010011100111: color_data = 12'b001110100111;
		16'b0000010011101000: color_data = 12'b001110100111;
		16'b0000010011101001: color_data = 12'b001110100111;
		16'b0000010011101010: color_data = 12'b001110100111;
		16'b0000010011101011: color_data = 12'b001110100111;
		16'b0000010011101100: color_data = 12'b001110100111;
		16'b0000010011101101: color_data = 12'b001110100111;
		16'b0000010011101110: color_data = 12'b001110100111;
		16'b0000010011101111: color_data = 12'b001110100111;
		16'b0000010011111100: color_data = 12'b001110100111;
		16'b0000010011111101: color_data = 12'b001110100111;
		16'b0000010011111110: color_data = 12'b001110100111;
		16'b0000010011111111: color_data = 12'b001110100111;
		16'b0000010100000000: color_data = 12'b001110100111;
		16'b0000010100000001: color_data = 12'b001110100111;
		16'b0000010100000010: color_data = 12'b001110100111;
		16'b0000010100000011: color_data = 12'b001110100111;
		16'b0000010100000100: color_data = 12'b001110100111;
		16'b0000010100000101: color_data = 12'b001110100111;
		16'b0000010100000110: color_data = 12'b001110100111;
		16'b0000010100000111: color_data = 12'b001110100111;
		16'b0000010100001000: color_data = 12'b001110100111;
		16'b0000010100001001: color_data = 12'b001110100111;
		16'b0000010100001010: color_data = 12'b001110100111;
		16'b0000010100001011: color_data = 12'b001110100111;
		16'b0000010100001100: color_data = 12'b001110100111;
		16'b0000010100001101: color_data = 12'b001110100111;
		16'b0000010100001110: color_data = 12'b001110100111;
		16'b0000010100001111: color_data = 12'b001110100111;
		16'b0000010100010000: color_data = 12'b001110100111;
		16'b0000010100010001: color_data = 12'b001110100111;
		16'b0000010100010010: color_data = 12'b001110100111;
		16'b0000010100010011: color_data = 12'b001110100111;
		16'b0000010100010100: color_data = 12'b001110100111;
		16'b0000010100010101: color_data = 12'b001110100111;
		16'b0000010100010110: color_data = 12'b001110100111;
		16'b0000010100010111: color_data = 12'b001110100111;
		16'b0000010100011000: color_data = 12'b001110100111;
		16'b0000010100011001: color_data = 12'b001110100111;
		16'b0000010100011010: color_data = 12'b001110100111;
		16'b0000010100011011: color_data = 12'b001110100111;
		16'b0000010100011100: color_data = 12'b001110100111;
		16'b0000010100011101: color_data = 12'b001110100111;
		16'b0000010100011110: color_data = 12'b001110100111;
		16'b0000010100011111: color_data = 12'b001110100111;
		16'b0000010100100000: color_data = 12'b001110100111;
		16'b0000010100101101: color_data = 12'b001110100111;
		16'b0000010100101110: color_data = 12'b001110100111;
		16'b0000010100101111: color_data = 12'b001110100111;
		16'b0000010100110000: color_data = 12'b001110100111;
		16'b0000010100110001: color_data = 12'b001110100111;
		16'b0000010100110010: color_data = 12'b001110100111;
		16'b0000010100110011: color_data = 12'b001110100111;
		16'b0000010100110100: color_data = 12'b001110100111;
		16'b0000010100110101: color_data = 12'b001110100111;
		16'b0000010100110110: color_data = 12'b001110100111;
		16'b0000010100110111: color_data = 12'b001110100111;
		16'b0000010100111000: color_data = 12'b001110100111;
		16'b0000010100111001: color_data = 12'b001110100111;
		16'b0000010100111010: color_data = 12'b001110100111;
		16'b0000010100111011: color_data = 12'b001110100111;
		16'b0000010100111100: color_data = 12'b001110100111;
		16'b0000010100111101: color_data = 12'b001110100111;
		16'b0000010100111110: color_data = 12'b001110100111;
		16'b0000010100111111: color_data = 12'b001110100111;
		16'b0000010101000000: color_data = 12'b001110100111;
		16'b0000010101000001: color_data = 12'b001110100111;
		16'b0000010101000010: color_data = 12'b001110100111;
		16'b0000010101000011: color_data = 12'b001110100111;
		16'b0000010101000100: color_data = 12'b001110100111;
		16'b0000010101100100: color_data = 12'b001110100111;
		16'b0000010101100101: color_data = 12'b001110100111;
		16'b0000010101100110: color_data = 12'b001110100111;
		16'b0000010101100111: color_data = 12'b001110100111;
		16'b0000010101101000: color_data = 12'b001110100111;
		16'b0000010101101001: color_data = 12'b001110100111;
		16'b0000010101101010: color_data = 12'b001110100111;
		16'b0000010101101011: color_data = 12'b001110100111;
		16'b0000010101101100: color_data = 12'b001110100111;
		16'b0000010101101101: color_data = 12'b001110100111;
		16'b0000010101101110: color_data = 12'b001110100111;
		16'b0000010101101111: color_data = 12'b001110100111;
		16'b0000010101110000: color_data = 12'b001110100111;
		16'b0000010101110001: color_data = 12'b001110100111;
		16'b0000010101110010: color_data = 12'b001110100111;
		16'b0000010101110011: color_data = 12'b001110100111;
		16'b0000010101110100: color_data = 12'b001110100111;
		16'b0000010101110101: color_data = 12'b001110100111;
		16'b0000010101110110: color_data = 12'b001110100111;
		16'b0000010101110111: color_data = 12'b001110100111;
		16'b0000010101111000: color_data = 12'b001110100111;
		16'b0000010101111001: color_data = 12'b001110100111;
		16'b0000010101111010: color_data = 12'b001110100111;
		16'b0000010101111011: color_data = 12'b001110100111;
		16'b0000011000001101: color_data = 12'b001110100111;
		16'b0000011000001110: color_data = 12'b001110100111;
		16'b0000011000001111: color_data = 12'b001110100111;
		16'b0000011000010000: color_data = 12'b001110100111;
		16'b0000011000010001: color_data = 12'b001110100111;
		16'b0000011000010010: color_data = 12'b001110100111;
		16'b0000011000010011: color_data = 12'b001110100111;
		16'b0000011000010100: color_data = 12'b001110100111;
		16'b0000011000010101: color_data = 12'b001110100111;
		16'b0000011000010110: color_data = 12'b001110100111;
		16'b0000011000010111: color_data = 12'b001110100111;
		16'b0000011000011000: color_data = 12'b001110100111;
		16'b0000011000011001: color_data = 12'b001110100111;
		16'b0000011000011010: color_data = 12'b001110100111;
		16'b0000011000011011: color_data = 12'b001110100111;
		16'b0000011000011100: color_data = 12'b001110100111;
		16'b0000011000011101: color_data = 12'b001110100111;
		16'b0000011000011110: color_data = 12'b001110100111;
		16'b0000011000011111: color_data = 12'b001110100111;
		16'b0000011000100000: color_data = 12'b001110100111;
		16'b0000011000100001: color_data = 12'b001110100111;
		16'b0000011000100010: color_data = 12'b001110100111;
		16'b0000011000100011: color_data = 12'b001110100111;
		16'b0000011000100100: color_data = 12'b001110100111;
		16'b0000011000101011: color_data = 12'b001110100111;
		16'b0000011000101100: color_data = 12'b001110100111;
		16'b0000011000101101: color_data = 12'b001110100111;
		16'b0000011000101110: color_data = 12'b001110100111;
		16'b0000011000101111: color_data = 12'b001110100111;
		16'b0000011000110000: color_data = 12'b001110100111;
		16'b0000011000110001: color_data = 12'b001110100111;
		16'b0000011000110010: color_data = 12'b001110100111;
		16'b0000011000110011: color_data = 12'b001110100111;
		16'b0000011000110100: color_data = 12'b001110100111;
		16'b0000011000110101: color_data = 12'b001110100111;
		16'b0000011000110110: color_data = 12'b001110100111;
		16'b0000011000110111: color_data = 12'b001110100111;
		16'b0000011001000100: color_data = 12'b001110100111;
		16'b0000011001000101: color_data = 12'b001110100111;
		16'b0000011001000110: color_data = 12'b001110100111;
		16'b0000011001000111: color_data = 12'b001110100111;
		16'b0000011001001000: color_data = 12'b001110100111;
		16'b0000011001001001: color_data = 12'b001110100111;
		16'b0000011001001010: color_data = 12'b001110100111;
		16'b0000011001001011: color_data = 12'b001110100111;
		16'b0000011001001100: color_data = 12'b001110100111;
		16'b0000011001001101: color_data = 12'b001110100111;
		16'b0000011001001110: color_data = 12'b001110100111;
		16'b0000011001001111: color_data = 12'b001110100111;
		16'b0000011001010110: color_data = 12'b001110100111;
		16'b0000011001010111: color_data = 12'b001110100111;
		16'b0000011001011000: color_data = 12'b001110100111;
		16'b0000011001011001: color_data = 12'b001110100111;
		16'b0000011001011010: color_data = 12'b001110100111;
		16'b0000011001011011: color_data = 12'b001110100111;
		16'b0000011001011100: color_data = 12'b001110100111;
		16'b0000011001011101: color_data = 12'b001110100111;
		16'b0000011001011110: color_data = 12'b001110100111;
		16'b0000011001011111: color_data = 12'b001110100111;
		16'b0000011001100000: color_data = 12'b001110100111;
		16'b0000011001100001: color_data = 12'b001110100111;
		16'b0000011001100010: color_data = 12'b001110100111;
		16'b0000011001100011: color_data = 12'b001110100111;
		16'b0000011001100100: color_data = 12'b001110100111;
		16'b0000011001100101: color_data = 12'b001110100111;
		16'b0000011001100110: color_data = 12'b001110100111;
		16'b0000011001100111: color_data = 12'b001110100111;
		16'b0000011001101000: color_data = 12'b001110100111;
		16'b0000011001101001: color_data = 12'b001110100111;
		16'b0000011001101010: color_data = 12'b001110100111;
		16'b0000011001101011: color_data = 12'b001110100111;
		16'b0000011001101100: color_data = 12'b001110100111;
		16'b0000011001101101: color_data = 12'b001110100111;
		16'b0000011001101110: color_data = 12'b001110100111;
		16'b0000011001110101: color_data = 12'b001110100111;
		16'b0000011001110110: color_data = 12'b001110100111;
		16'b0000011001110111: color_data = 12'b001110100111;
		16'b0000011001111000: color_data = 12'b001110100111;
		16'b0000011001111001: color_data = 12'b001110100111;
		16'b0000011001111010: color_data = 12'b001110100111;
		16'b0000011001111011: color_data = 12'b001110100111;
		16'b0000011001111100: color_data = 12'b001110100111;
		16'b0000011001111101: color_data = 12'b001110100111;
		16'b0000011001111110: color_data = 12'b001110100111;
		16'b0000011001111111: color_data = 12'b001110100111;
		16'b0000011010000000: color_data = 12'b001110100111;
		16'b0000011010000001: color_data = 12'b001110100111;
		16'b0000011010000010: color_data = 12'b001110100111;
		16'b0000011010000011: color_data = 12'b001110100111;
		16'b0000011010000100: color_data = 12'b001110100111;
		16'b0000011010000101: color_data = 12'b001110100111;
		16'b0000011010000110: color_data = 12'b001110100111;
		16'b0000011010000111: color_data = 12'b001110100111;
		16'b0000011010001000: color_data = 12'b001110100111;
		16'b0000011010001001: color_data = 12'b001110100111;
		16'b0000011010001010: color_data = 12'b001110100111;
		16'b0000011010001011: color_data = 12'b001110100111;
		16'b0000011010001100: color_data = 12'b001110100111;
		16'b0000011010101100: color_data = 12'b001110100111;
		16'b0000011010101101: color_data = 12'b001110100111;
		16'b0000011010101110: color_data = 12'b001110100111;
		16'b0000011010101111: color_data = 12'b001110100111;
		16'b0000011010110000: color_data = 12'b001110100111;
		16'b0000011010110001: color_data = 12'b001110100111;
		16'b0000011010110010: color_data = 12'b001110100111;
		16'b0000011010110011: color_data = 12'b001110100111;
		16'b0000011010110100: color_data = 12'b001110100111;
		16'b0000011010110101: color_data = 12'b001110100111;
		16'b0000011010110110: color_data = 12'b001110100111;
		16'b0000011010110111: color_data = 12'b001110100111;
		16'b0000011010111000: color_data = 12'b001110100111;
		16'b0000011010111001: color_data = 12'b001110100111;
		16'b0000011010111010: color_data = 12'b001110100111;
		16'b0000011010111011: color_data = 12'b001110100111;
		16'b0000011010111100: color_data = 12'b001110100111;
		16'b0000011010111101: color_data = 12'b001110100111;
		16'b0000011010111110: color_data = 12'b001110100111;
		16'b0000011010111111: color_data = 12'b001110100111;
		16'b0000011011000000: color_data = 12'b001110100111;
		16'b0000011011000001: color_data = 12'b001110100111;
		16'b0000011011000010: color_data = 12'b001110100111;
		16'b0000011011000011: color_data = 12'b001110100111;
		16'b0000011011000100: color_data = 12'b001110100111;
		16'b0000011011001011: color_data = 12'b001110100111;
		16'b0000011011001100: color_data = 12'b001110100111;
		16'b0000011011001101: color_data = 12'b001110100111;
		16'b0000011011001110: color_data = 12'b001110100111;
		16'b0000011011001111: color_data = 12'b001110100111;
		16'b0000011011010000: color_data = 12'b001110100111;
		16'b0000011011010001: color_data = 12'b001110100111;
		16'b0000011011010010: color_data = 12'b001110100111;
		16'b0000011011010011: color_data = 12'b001110100111;
		16'b0000011011010100: color_data = 12'b001110100111;
		16'b0000011011010101: color_data = 12'b001110100111;
		16'b0000011011010110: color_data = 12'b001110100111;
		16'b0000011011010111: color_data = 12'b001110100111;
		16'b0000011011011000: color_data = 12'b001110100111;
		16'b0000011011011001: color_data = 12'b001110100111;
		16'b0000011011011010: color_data = 12'b001110100111;
		16'b0000011011011011: color_data = 12'b001110100111;
		16'b0000011011011100: color_data = 12'b001110100111;
		16'b0000011011011101: color_data = 12'b001110100111;
		16'b0000011011011110: color_data = 12'b001110100111;
		16'b0000011011011111: color_data = 12'b001110100111;
		16'b0000011011100000: color_data = 12'b001110100111;
		16'b0000011011100001: color_data = 12'b001110100111;
		16'b0000011011100010: color_data = 12'b001110100111;
		16'b0000011011100011: color_data = 12'b001110100111;
		16'b0000011011100100: color_data = 12'b001110100111;
		16'b0000011011100101: color_data = 12'b001110100111;
		16'b0000011011100110: color_data = 12'b001110100111;
		16'b0000011011100111: color_data = 12'b001110100111;
		16'b0000011011101000: color_data = 12'b001110100111;
		16'b0000011011101001: color_data = 12'b001110100111;
		16'b0000011011101010: color_data = 12'b001110100111;
		16'b0000011011101011: color_data = 12'b001110100111;
		16'b0000011011101100: color_data = 12'b001110100111;
		16'b0000011011101101: color_data = 12'b001110100111;
		16'b0000011011101110: color_data = 12'b001110100111;
		16'b0000011011101111: color_data = 12'b001110100111;
		16'b0000011011111100: color_data = 12'b001110100111;
		16'b0000011011111101: color_data = 12'b001110100111;
		16'b0000011011111110: color_data = 12'b001110100111;
		16'b0000011011111111: color_data = 12'b001110100111;
		16'b0000011100000000: color_data = 12'b001110100111;
		16'b0000011100000001: color_data = 12'b001110100111;
		16'b0000011100000010: color_data = 12'b001110100111;
		16'b0000011100000011: color_data = 12'b001110100111;
		16'b0000011100000100: color_data = 12'b001110100111;
		16'b0000011100000101: color_data = 12'b001110100111;
		16'b0000011100000110: color_data = 12'b001110100111;
		16'b0000011100000111: color_data = 12'b001110100111;
		16'b0000011100001000: color_data = 12'b001110100111;
		16'b0000011100001001: color_data = 12'b001110100111;
		16'b0000011100001010: color_data = 12'b001110100111;
		16'b0000011100001011: color_data = 12'b001110100111;
		16'b0000011100001100: color_data = 12'b001110100111;
		16'b0000011100001101: color_data = 12'b001110100111;
		16'b0000011100001110: color_data = 12'b001110100111;
		16'b0000011100001111: color_data = 12'b001110100111;
		16'b0000011100010000: color_data = 12'b001110100111;
		16'b0000011100010001: color_data = 12'b001110100111;
		16'b0000011100010010: color_data = 12'b001110100111;
		16'b0000011100010011: color_data = 12'b001110100111;
		16'b0000011100010100: color_data = 12'b001110100111;
		16'b0000011100010101: color_data = 12'b001110100111;
		16'b0000011100010110: color_data = 12'b001110100111;
		16'b0000011100010111: color_data = 12'b001110100111;
		16'b0000011100011000: color_data = 12'b001110100111;
		16'b0000011100011001: color_data = 12'b001110100111;
		16'b0000011100011010: color_data = 12'b001110100111;
		16'b0000011100011011: color_data = 12'b001110100111;
		16'b0000011100011100: color_data = 12'b001110100111;
		16'b0000011100011101: color_data = 12'b001110100111;
		16'b0000011100011110: color_data = 12'b001110100111;
		16'b0000011100011111: color_data = 12'b001110100111;
		16'b0000011100100000: color_data = 12'b001110100111;
		16'b0000011100101101: color_data = 12'b001110100111;
		16'b0000011100101110: color_data = 12'b001110100111;
		16'b0000011100101111: color_data = 12'b001110100111;
		16'b0000011100110000: color_data = 12'b001110100111;
		16'b0000011100110001: color_data = 12'b001110100111;
		16'b0000011100110010: color_data = 12'b001110100111;
		16'b0000011100110011: color_data = 12'b001110100111;
		16'b0000011100110100: color_data = 12'b001110100111;
		16'b0000011100110101: color_data = 12'b001110100111;
		16'b0000011100110110: color_data = 12'b001110100111;
		16'b0000011100110111: color_data = 12'b001110100111;
		16'b0000011100111000: color_data = 12'b001110100111;
		16'b0000011100111001: color_data = 12'b001110100111;
		16'b0000011100111010: color_data = 12'b001110100111;
		16'b0000011100111011: color_data = 12'b001110100111;
		16'b0000011100111100: color_data = 12'b001110100111;
		16'b0000011100111101: color_data = 12'b001110100111;
		16'b0000011100111110: color_data = 12'b001110100111;
		16'b0000011100111111: color_data = 12'b001110100111;
		16'b0000011101000000: color_data = 12'b001110100111;
		16'b0000011101000001: color_data = 12'b001110100111;
		16'b0000011101000010: color_data = 12'b001110100111;
		16'b0000011101000011: color_data = 12'b001110100111;
		16'b0000011101000100: color_data = 12'b001110100111;
		16'b0000011101100100: color_data = 12'b001110100111;
		16'b0000011101100101: color_data = 12'b001110100111;
		16'b0000011101100110: color_data = 12'b001110100111;
		16'b0000011101100111: color_data = 12'b001110100111;
		16'b0000011101101000: color_data = 12'b001110100111;
		16'b0000011101101001: color_data = 12'b001110100111;
		16'b0000011101101010: color_data = 12'b001110100111;
		16'b0000011101101011: color_data = 12'b001110100111;
		16'b0000011101101100: color_data = 12'b001110100111;
		16'b0000011101101101: color_data = 12'b001110100111;
		16'b0000011101101110: color_data = 12'b001110100111;
		16'b0000011101101111: color_data = 12'b001110100111;
		16'b0000011101110000: color_data = 12'b001110100111;
		16'b0000011101110001: color_data = 12'b001110100111;
		16'b0000011101110010: color_data = 12'b001110100111;
		16'b0000011101110011: color_data = 12'b001110100111;
		16'b0000011101110100: color_data = 12'b001110100111;
		16'b0000011101110101: color_data = 12'b001110100111;
		16'b0000011101110110: color_data = 12'b001110100111;
		16'b0000011101110111: color_data = 12'b001110100111;
		16'b0000011101111000: color_data = 12'b001110100111;
		16'b0000011101111001: color_data = 12'b001110100111;
		16'b0000011101111010: color_data = 12'b001110100111;
		16'b0000011101111011: color_data = 12'b001110100111;
		16'b0000100000001101: color_data = 12'b001110100111;
		16'b0000100000001110: color_data = 12'b001110100111;
		16'b0000100000001111: color_data = 12'b001110100111;
		16'b0000100000010000: color_data = 12'b001110100111;
		16'b0000100000010001: color_data = 12'b001110100111;
		16'b0000100000010010: color_data = 12'b001110100111;
		16'b0000100000010011: color_data = 12'b001110100111;
		16'b0000100000010100: color_data = 12'b001110100111;
		16'b0000100000010101: color_data = 12'b001110100111;
		16'b0000100000010110: color_data = 12'b001110100111;
		16'b0000100000010111: color_data = 12'b001110100111;
		16'b0000100000011000: color_data = 12'b001110100111;
		16'b0000100000011001: color_data = 12'b001110100111;
		16'b0000100000011010: color_data = 12'b001110100111;
		16'b0000100000011011: color_data = 12'b001110100111;
		16'b0000100000011100: color_data = 12'b001110100111;
		16'b0000100000011101: color_data = 12'b001110100111;
		16'b0000100000011110: color_data = 12'b001110100111;
		16'b0000100000011111: color_data = 12'b001110100111;
		16'b0000100000100000: color_data = 12'b001110100111;
		16'b0000100000100001: color_data = 12'b001110100111;
		16'b0000100000100010: color_data = 12'b001110100111;
		16'b0000100000100011: color_data = 12'b001110100111;
		16'b0000100000100100: color_data = 12'b001110100111;
		16'b0000100000101011: color_data = 12'b001110100111;
		16'b0000100000101100: color_data = 12'b001110100111;
		16'b0000100000101101: color_data = 12'b001110100111;
		16'b0000100000101110: color_data = 12'b001110100111;
		16'b0000100000101111: color_data = 12'b001110100111;
		16'b0000100000110000: color_data = 12'b001110100111;
		16'b0000100000110001: color_data = 12'b001110100111;
		16'b0000100000110010: color_data = 12'b001110100111;
		16'b0000100000110011: color_data = 12'b001110100111;
		16'b0000100000110100: color_data = 12'b001110100111;
		16'b0000100000110101: color_data = 12'b001110100111;
		16'b0000100000110110: color_data = 12'b001110100111;
		16'b0000100000110111: color_data = 12'b001110100111;
		16'b0000100001000100: color_data = 12'b001110100111;
		16'b0000100001000101: color_data = 12'b001110100111;
		16'b0000100001000110: color_data = 12'b001110100111;
		16'b0000100001000111: color_data = 12'b001110100111;
		16'b0000100001001000: color_data = 12'b001110100111;
		16'b0000100001001001: color_data = 12'b001110100111;
		16'b0000100001001010: color_data = 12'b001110100111;
		16'b0000100001001011: color_data = 12'b001110100111;
		16'b0000100001001100: color_data = 12'b001110100111;
		16'b0000100001001101: color_data = 12'b001110100111;
		16'b0000100001001110: color_data = 12'b001110100111;
		16'b0000100001001111: color_data = 12'b001110100111;
		16'b0000100001010110: color_data = 12'b001110100111;
		16'b0000100001010111: color_data = 12'b001110100111;
		16'b0000100001011000: color_data = 12'b001110100111;
		16'b0000100001011001: color_data = 12'b001110100111;
		16'b0000100001011010: color_data = 12'b001110100111;
		16'b0000100001011011: color_data = 12'b001110100111;
		16'b0000100001011100: color_data = 12'b001110100111;
		16'b0000100001011101: color_data = 12'b001110100111;
		16'b0000100001011110: color_data = 12'b001110100111;
		16'b0000100001011111: color_data = 12'b001110100111;
		16'b0000100001100000: color_data = 12'b001110100111;
		16'b0000100001100001: color_data = 12'b001110100111;
		16'b0000100001100010: color_data = 12'b001110100111;
		16'b0000100001100011: color_data = 12'b001110100111;
		16'b0000100001100100: color_data = 12'b001110100111;
		16'b0000100001100101: color_data = 12'b001110100111;
		16'b0000100001100110: color_data = 12'b001110100111;
		16'b0000100001100111: color_data = 12'b001110100111;
		16'b0000100001101000: color_data = 12'b001110100111;
		16'b0000100001101001: color_data = 12'b001110100111;
		16'b0000100001101010: color_data = 12'b001110100111;
		16'b0000100001101011: color_data = 12'b001110100111;
		16'b0000100001101100: color_data = 12'b001110100111;
		16'b0000100001101101: color_data = 12'b001110100111;
		16'b0000100001101110: color_data = 12'b001110100111;
		16'b0000100001110101: color_data = 12'b001110100111;
		16'b0000100001110110: color_data = 12'b001110100111;
		16'b0000100001110111: color_data = 12'b001110100111;
		16'b0000100001111000: color_data = 12'b001110100111;
		16'b0000100001111001: color_data = 12'b001110100111;
		16'b0000100001111010: color_data = 12'b001110100111;
		16'b0000100001111011: color_data = 12'b001110100111;
		16'b0000100001111100: color_data = 12'b001110100111;
		16'b0000100001111101: color_data = 12'b001110100111;
		16'b0000100001111110: color_data = 12'b001110100111;
		16'b0000100001111111: color_data = 12'b001110100111;
		16'b0000100010000000: color_data = 12'b001110100111;
		16'b0000100010000001: color_data = 12'b001110100111;
		16'b0000100010000010: color_data = 12'b001110100111;
		16'b0000100010000011: color_data = 12'b001110100111;
		16'b0000100010000100: color_data = 12'b001110100111;
		16'b0000100010000101: color_data = 12'b001110100111;
		16'b0000100010000110: color_data = 12'b001110100111;
		16'b0000100010000111: color_data = 12'b001110100111;
		16'b0000100010001000: color_data = 12'b001110100111;
		16'b0000100010001001: color_data = 12'b001110100111;
		16'b0000100010001010: color_data = 12'b001110100111;
		16'b0000100010001011: color_data = 12'b001110100111;
		16'b0000100010001100: color_data = 12'b001110100111;
		16'b0000100010101100: color_data = 12'b001110100111;
		16'b0000100010101101: color_data = 12'b001110100111;
		16'b0000100010101110: color_data = 12'b001110100111;
		16'b0000100010101111: color_data = 12'b001110100111;
		16'b0000100010110000: color_data = 12'b001110100111;
		16'b0000100010110001: color_data = 12'b001110100111;
		16'b0000100010110010: color_data = 12'b001110100111;
		16'b0000100010110011: color_data = 12'b001110100111;
		16'b0000100010110100: color_data = 12'b001110100111;
		16'b0000100010110101: color_data = 12'b001110100111;
		16'b0000100010110110: color_data = 12'b001110100111;
		16'b0000100010110111: color_data = 12'b001110100111;
		16'b0000100010111000: color_data = 12'b001110100111;
		16'b0000100010111001: color_data = 12'b001110100111;
		16'b0000100010111010: color_data = 12'b001110100111;
		16'b0000100010111011: color_data = 12'b001110100111;
		16'b0000100010111100: color_data = 12'b001110100111;
		16'b0000100010111101: color_data = 12'b001110100111;
		16'b0000100010111110: color_data = 12'b001110100111;
		16'b0000100010111111: color_data = 12'b001110100111;
		16'b0000100011000000: color_data = 12'b001110100111;
		16'b0000100011000001: color_data = 12'b001110100111;
		16'b0000100011000010: color_data = 12'b001110100111;
		16'b0000100011000011: color_data = 12'b001110100111;
		16'b0000100011000100: color_data = 12'b001110100111;
		16'b0000100011001011: color_data = 12'b001110100111;
		16'b0000100011001100: color_data = 12'b001110100111;
		16'b0000100011001101: color_data = 12'b001110100111;
		16'b0000100011001110: color_data = 12'b001110100111;
		16'b0000100011001111: color_data = 12'b001110100111;
		16'b0000100011010000: color_data = 12'b001110100111;
		16'b0000100011010001: color_data = 12'b001110100111;
		16'b0000100011010010: color_data = 12'b001110100111;
		16'b0000100011010011: color_data = 12'b001110100111;
		16'b0000100011010100: color_data = 12'b001110100111;
		16'b0000100011010101: color_data = 12'b001110100111;
		16'b0000100011010110: color_data = 12'b001110100111;
		16'b0000100011010111: color_data = 12'b001110100111;
		16'b0000100011011000: color_data = 12'b001110100111;
		16'b0000100011011001: color_data = 12'b001110100111;
		16'b0000100011011010: color_data = 12'b001110100111;
		16'b0000100011011011: color_data = 12'b001110100111;
		16'b0000100011011100: color_data = 12'b001110100111;
		16'b0000100011011101: color_data = 12'b001110100111;
		16'b0000100011011110: color_data = 12'b001110100111;
		16'b0000100011011111: color_data = 12'b001110100111;
		16'b0000100011100000: color_data = 12'b001110100111;
		16'b0000100011100001: color_data = 12'b001110100111;
		16'b0000100011100010: color_data = 12'b001110100111;
		16'b0000100011100011: color_data = 12'b001110100111;
		16'b0000100011100100: color_data = 12'b001110100111;
		16'b0000100011100101: color_data = 12'b001110100111;
		16'b0000100011100110: color_data = 12'b001110100111;
		16'b0000100011100111: color_data = 12'b001110100111;
		16'b0000100011101000: color_data = 12'b001110100111;
		16'b0000100011101001: color_data = 12'b001110100111;
		16'b0000100011101010: color_data = 12'b001110100111;
		16'b0000100011101011: color_data = 12'b001110100111;
		16'b0000100011101100: color_data = 12'b001110100111;
		16'b0000100011101101: color_data = 12'b001110100111;
		16'b0000100011101110: color_data = 12'b001110100111;
		16'b0000100011101111: color_data = 12'b001110100111;
		16'b0000100011111100: color_data = 12'b001110100111;
		16'b0000100011111101: color_data = 12'b001110100111;
		16'b0000100011111110: color_data = 12'b001110100111;
		16'b0000100011111111: color_data = 12'b001110100111;
		16'b0000100100000000: color_data = 12'b001110100111;
		16'b0000100100000001: color_data = 12'b001110100111;
		16'b0000100100000010: color_data = 12'b001110100111;
		16'b0000100100000011: color_data = 12'b001110100111;
		16'b0000100100000100: color_data = 12'b001110100111;
		16'b0000100100000101: color_data = 12'b001110100111;
		16'b0000100100000110: color_data = 12'b001110100111;
		16'b0000100100000111: color_data = 12'b001110100111;
		16'b0000100100001000: color_data = 12'b001110100111;
		16'b0000100100001001: color_data = 12'b001110100111;
		16'b0000100100001010: color_data = 12'b001110100111;
		16'b0000100100001011: color_data = 12'b001110100111;
		16'b0000100100001100: color_data = 12'b001110100111;
		16'b0000100100001101: color_data = 12'b001110100111;
		16'b0000100100001110: color_data = 12'b001110100111;
		16'b0000100100001111: color_data = 12'b001110100111;
		16'b0000100100010000: color_data = 12'b001110100111;
		16'b0000100100010001: color_data = 12'b001110100111;
		16'b0000100100010010: color_data = 12'b001110100111;
		16'b0000100100010011: color_data = 12'b001110100111;
		16'b0000100100010100: color_data = 12'b001110100111;
		16'b0000100100010101: color_data = 12'b001110100111;
		16'b0000100100010110: color_data = 12'b001110100111;
		16'b0000100100010111: color_data = 12'b001110100111;
		16'b0000100100011000: color_data = 12'b001110100111;
		16'b0000100100011001: color_data = 12'b001110100111;
		16'b0000100100011010: color_data = 12'b001110100111;
		16'b0000100100011011: color_data = 12'b001110100111;
		16'b0000100100011100: color_data = 12'b001110100111;
		16'b0000100100011101: color_data = 12'b001110100111;
		16'b0000100100011110: color_data = 12'b001110100111;
		16'b0000100100011111: color_data = 12'b001110100111;
		16'b0000100100100000: color_data = 12'b001110100111;
		16'b0000100100101101: color_data = 12'b001110100111;
		16'b0000100100101110: color_data = 12'b001110100111;
		16'b0000100100101111: color_data = 12'b001110100111;
		16'b0000100100110000: color_data = 12'b001110100111;
		16'b0000100100110001: color_data = 12'b001110100111;
		16'b0000100100110010: color_data = 12'b001110100111;
		16'b0000100100110011: color_data = 12'b001110100111;
		16'b0000100100110100: color_data = 12'b001110100111;
		16'b0000100100110101: color_data = 12'b001110100111;
		16'b0000100100110110: color_data = 12'b001110100111;
		16'b0000100100110111: color_data = 12'b001110100111;
		16'b0000100100111000: color_data = 12'b001110100111;
		16'b0000100100111001: color_data = 12'b001110100111;
		16'b0000100100111010: color_data = 12'b001110100111;
		16'b0000100100111011: color_data = 12'b001110100111;
		16'b0000100100111100: color_data = 12'b001110100111;
		16'b0000100100111101: color_data = 12'b001110100111;
		16'b0000100100111110: color_data = 12'b001110100111;
		16'b0000100100111111: color_data = 12'b001110100111;
		16'b0000100101000000: color_data = 12'b001110100111;
		16'b0000100101000001: color_data = 12'b001110100111;
		16'b0000100101000010: color_data = 12'b001110100111;
		16'b0000100101000011: color_data = 12'b001110100111;
		16'b0000100101000100: color_data = 12'b001110100111;
		16'b0000100101100100: color_data = 12'b001110100111;
		16'b0000100101100101: color_data = 12'b001110100111;
		16'b0000100101100110: color_data = 12'b001110100111;
		16'b0000100101100111: color_data = 12'b001110100111;
		16'b0000100101101000: color_data = 12'b001110100111;
		16'b0000100101101001: color_data = 12'b001110100111;
		16'b0000100101101010: color_data = 12'b001110100111;
		16'b0000100101101011: color_data = 12'b001110100111;
		16'b0000100101101100: color_data = 12'b001110100111;
		16'b0000100101101101: color_data = 12'b001110100111;
		16'b0000100101101110: color_data = 12'b001110100111;
		16'b0000100101101111: color_data = 12'b001110100111;
		16'b0000100101110000: color_data = 12'b001110100111;
		16'b0000100101110001: color_data = 12'b001110100111;
		16'b0000100101110010: color_data = 12'b001110100111;
		16'b0000100101110011: color_data = 12'b001110100111;
		16'b0000100101110100: color_data = 12'b001110100111;
		16'b0000100101110101: color_data = 12'b001110100111;
		16'b0000100101110110: color_data = 12'b001110100111;
		16'b0000100101110111: color_data = 12'b001110100111;
		16'b0000100101111000: color_data = 12'b001110100111;
		16'b0000100101111001: color_data = 12'b001110100111;
		16'b0000100101111010: color_data = 12'b001110100111;
		16'b0000100101111011: color_data = 12'b001110100111;
		16'b0000101000001101: color_data = 12'b001110100111;
		16'b0000101000001110: color_data = 12'b001110100111;
		16'b0000101000001111: color_data = 12'b001110100111;
		16'b0000101000010000: color_data = 12'b001110100111;
		16'b0000101000010001: color_data = 12'b001110100111;
		16'b0000101000010010: color_data = 12'b001110100111;
		16'b0000101000010011: color_data = 12'b001110100111;
		16'b0000101000010100: color_data = 12'b001110100111;
		16'b0000101000010101: color_data = 12'b001110100111;
		16'b0000101000010110: color_data = 12'b001110100111;
		16'b0000101000010111: color_data = 12'b001110100111;
		16'b0000101000011000: color_data = 12'b001110100111;
		16'b0000101000011001: color_data = 12'b001110100111;
		16'b0000101000011010: color_data = 12'b001110100111;
		16'b0000101000011011: color_data = 12'b001110100111;
		16'b0000101000011100: color_data = 12'b001110100111;
		16'b0000101000011101: color_data = 12'b001110100111;
		16'b0000101000011110: color_data = 12'b001110100111;
		16'b0000101000011111: color_data = 12'b001110100111;
		16'b0000101000100000: color_data = 12'b001110100111;
		16'b0000101000100001: color_data = 12'b001110100111;
		16'b0000101000100010: color_data = 12'b001110100111;
		16'b0000101000100011: color_data = 12'b001110100111;
		16'b0000101000100100: color_data = 12'b001110100111;
		16'b0000101000101011: color_data = 12'b001110100111;
		16'b0000101000101100: color_data = 12'b001110100111;
		16'b0000101000101101: color_data = 12'b001110100111;
		16'b0000101000101110: color_data = 12'b001110100111;
		16'b0000101000101111: color_data = 12'b001110100111;
		16'b0000101000110000: color_data = 12'b001110100111;
		16'b0000101000110001: color_data = 12'b001110100111;
		16'b0000101000110010: color_data = 12'b001110100111;
		16'b0000101000110011: color_data = 12'b001110100111;
		16'b0000101000110100: color_data = 12'b001110100111;
		16'b0000101000110101: color_data = 12'b001110100111;
		16'b0000101000110110: color_data = 12'b001110100111;
		16'b0000101000110111: color_data = 12'b001110100111;
		16'b0000101001000100: color_data = 12'b001110100111;
		16'b0000101001000101: color_data = 12'b001110100111;
		16'b0000101001000110: color_data = 12'b001110100111;
		16'b0000101001000111: color_data = 12'b001110100111;
		16'b0000101001001000: color_data = 12'b001110100111;
		16'b0000101001001001: color_data = 12'b001110100111;
		16'b0000101001001010: color_data = 12'b001110100111;
		16'b0000101001001011: color_data = 12'b001110100111;
		16'b0000101001001100: color_data = 12'b001110100111;
		16'b0000101001001101: color_data = 12'b001110100111;
		16'b0000101001001110: color_data = 12'b001110100111;
		16'b0000101001001111: color_data = 12'b001110100111;
		16'b0000101001010110: color_data = 12'b001110100111;
		16'b0000101001010111: color_data = 12'b001110100111;
		16'b0000101001011000: color_data = 12'b001110100111;
		16'b0000101001011001: color_data = 12'b001110100111;
		16'b0000101001011010: color_data = 12'b001110100111;
		16'b0000101001011011: color_data = 12'b001110100111;
		16'b0000101001011100: color_data = 12'b001110100111;
		16'b0000101001011101: color_data = 12'b001110100111;
		16'b0000101001011110: color_data = 12'b001110100111;
		16'b0000101001011111: color_data = 12'b001110100111;
		16'b0000101001100000: color_data = 12'b001110100111;
		16'b0000101001100001: color_data = 12'b001110100111;
		16'b0000101001100010: color_data = 12'b001110100111;
		16'b0000101001100011: color_data = 12'b001110100111;
		16'b0000101001100100: color_data = 12'b001110100111;
		16'b0000101001100101: color_data = 12'b001110100111;
		16'b0000101001100110: color_data = 12'b001110100111;
		16'b0000101001100111: color_data = 12'b001110100111;
		16'b0000101001101000: color_data = 12'b001110100111;
		16'b0000101001101001: color_data = 12'b001110100111;
		16'b0000101001101010: color_data = 12'b001110100111;
		16'b0000101001101011: color_data = 12'b001110100111;
		16'b0000101001101100: color_data = 12'b001110100111;
		16'b0000101001101101: color_data = 12'b001110100111;
		16'b0000101001101110: color_data = 12'b001110100111;
		16'b0000101001110101: color_data = 12'b001110100111;
		16'b0000101001110110: color_data = 12'b001110100111;
		16'b0000101001110111: color_data = 12'b001110100111;
		16'b0000101001111000: color_data = 12'b001110100111;
		16'b0000101001111001: color_data = 12'b001110100111;
		16'b0000101001111010: color_data = 12'b001110100111;
		16'b0000101001111011: color_data = 12'b001110100111;
		16'b0000101001111100: color_data = 12'b001110100111;
		16'b0000101001111101: color_data = 12'b001110100111;
		16'b0000101001111110: color_data = 12'b001110100111;
		16'b0000101001111111: color_data = 12'b001110100111;
		16'b0000101010000000: color_data = 12'b001110100111;
		16'b0000101010000001: color_data = 12'b001110100111;
		16'b0000101010000010: color_data = 12'b001110100111;
		16'b0000101010000011: color_data = 12'b001110100111;
		16'b0000101010000100: color_data = 12'b001110100111;
		16'b0000101010000101: color_data = 12'b001110100111;
		16'b0000101010000110: color_data = 12'b001110100111;
		16'b0000101010000111: color_data = 12'b001110100111;
		16'b0000101010001000: color_data = 12'b001110100111;
		16'b0000101010001001: color_data = 12'b001110100111;
		16'b0000101010001010: color_data = 12'b001110100111;
		16'b0000101010001011: color_data = 12'b001110100111;
		16'b0000101010001100: color_data = 12'b001110100111;
		16'b0000101010101100: color_data = 12'b001110100111;
		16'b0000101010101101: color_data = 12'b001110100111;
		16'b0000101010101110: color_data = 12'b001110100111;
		16'b0000101010101111: color_data = 12'b001110100111;
		16'b0000101010110000: color_data = 12'b001110100111;
		16'b0000101010110001: color_data = 12'b001110100111;
		16'b0000101010110010: color_data = 12'b001110100111;
		16'b0000101010110011: color_data = 12'b001110100111;
		16'b0000101010110100: color_data = 12'b001110100111;
		16'b0000101010110101: color_data = 12'b001110100111;
		16'b0000101010110110: color_data = 12'b001110100111;
		16'b0000101010110111: color_data = 12'b001110100111;
		16'b0000101010111000: color_data = 12'b001110100111;
		16'b0000101010111001: color_data = 12'b001110100111;
		16'b0000101010111010: color_data = 12'b001110100111;
		16'b0000101010111011: color_data = 12'b001110100111;
		16'b0000101010111100: color_data = 12'b001110100111;
		16'b0000101010111101: color_data = 12'b001110100111;
		16'b0000101010111110: color_data = 12'b001110100111;
		16'b0000101010111111: color_data = 12'b001110100111;
		16'b0000101011000000: color_data = 12'b001110100111;
		16'b0000101011000001: color_data = 12'b001110100111;
		16'b0000101011000010: color_data = 12'b001110100111;
		16'b0000101011000011: color_data = 12'b001110100111;
		16'b0000101011000100: color_data = 12'b001110100111;
		16'b0000101011001011: color_data = 12'b001110100111;
		16'b0000101011001100: color_data = 12'b001110100111;
		16'b0000101011001101: color_data = 12'b001110100111;
		16'b0000101011001110: color_data = 12'b001110100111;
		16'b0000101011001111: color_data = 12'b001110100111;
		16'b0000101011010000: color_data = 12'b001110100111;
		16'b0000101011010001: color_data = 12'b001110100111;
		16'b0000101011010010: color_data = 12'b001110100111;
		16'b0000101011010011: color_data = 12'b001110100111;
		16'b0000101011010100: color_data = 12'b001110100111;
		16'b0000101011010101: color_data = 12'b001110100111;
		16'b0000101011010110: color_data = 12'b001110100111;
		16'b0000101011010111: color_data = 12'b001110100111;
		16'b0000101011011000: color_data = 12'b001110100111;
		16'b0000101011011001: color_data = 12'b001110100111;
		16'b0000101011011010: color_data = 12'b001110100111;
		16'b0000101011011011: color_data = 12'b001110100111;
		16'b0000101011011100: color_data = 12'b001110100111;
		16'b0000101011011101: color_data = 12'b001110100111;
		16'b0000101011011110: color_data = 12'b001110100111;
		16'b0000101011011111: color_data = 12'b001110100111;
		16'b0000101011100000: color_data = 12'b001110100111;
		16'b0000101011100001: color_data = 12'b001110100111;
		16'b0000101011100010: color_data = 12'b001110100111;
		16'b0000101011100011: color_data = 12'b001110100111;
		16'b0000101011100100: color_data = 12'b001110100111;
		16'b0000101011100101: color_data = 12'b001110100111;
		16'b0000101011100110: color_data = 12'b001110100111;
		16'b0000101011100111: color_data = 12'b001110100111;
		16'b0000101011101000: color_data = 12'b001110100111;
		16'b0000101011101001: color_data = 12'b001110100111;
		16'b0000101011101010: color_data = 12'b001110100111;
		16'b0000101011101011: color_data = 12'b001110100111;
		16'b0000101011101100: color_data = 12'b001110100111;
		16'b0000101011101101: color_data = 12'b001110100111;
		16'b0000101011101110: color_data = 12'b001110100111;
		16'b0000101011101111: color_data = 12'b001110100111;
		16'b0000101011111100: color_data = 12'b001110100111;
		16'b0000101011111101: color_data = 12'b001110100111;
		16'b0000101011111110: color_data = 12'b001110100111;
		16'b0000101011111111: color_data = 12'b001110100111;
		16'b0000101100000000: color_data = 12'b001110100111;
		16'b0000101100000001: color_data = 12'b001110100111;
		16'b0000101100000010: color_data = 12'b001110100111;
		16'b0000101100000011: color_data = 12'b001110100111;
		16'b0000101100000100: color_data = 12'b001110100111;
		16'b0000101100000101: color_data = 12'b001110100111;
		16'b0000101100000110: color_data = 12'b001110100111;
		16'b0000101100000111: color_data = 12'b001110100111;
		16'b0000101100001000: color_data = 12'b001110100111;
		16'b0000101100001001: color_data = 12'b001110100111;
		16'b0000101100001010: color_data = 12'b001110100111;
		16'b0000101100001011: color_data = 12'b001110100111;
		16'b0000101100001100: color_data = 12'b001110100111;
		16'b0000101100001101: color_data = 12'b001110100111;
		16'b0000101100001110: color_data = 12'b001110100111;
		16'b0000101100001111: color_data = 12'b001110100111;
		16'b0000101100010000: color_data = 12'b001110100111;
		16'b0000101100010001: color_data = 12'b001110100111;
		16'b0000101100010010: color_data = 12'b001110100111;
		16'b0000101100010011: color_data = 12'b001110100111;
		16'b0000101100010100: color_data = 12'b001110100111;
		16'b0000101100010101: color_data = 12'b001110100111;
		16'b0000101100010110: color_data = 12'b001110100111;
		16'b0000101100010111: color_data = 12'b001110100111;
		16'b0000101100011000: color_data = 12'b001110100111;
		16'b0000101100011001: color_data = 12'b001110100111;
		16'b0000101100011010: color_data = 12'b001110100111;
		16'b0000101100011011: color_data = 12'b001110100111;
		16'b0000101100011100: color_data = 12'b001110100111;
		16'b0000101100011101: color_data = 12'b001110100111;
		16'b0000101100011110: color_data = 12'b001110100111;
		16'b0000101100011111: color_data = 12'b001110100111;
		16'b0000101100100000: color_data = 12'b001110100111;
		16'b0000101100101101: color_data = 12'b001110100111;
		16'b0000101100101110: color_data = 12'b001110100111;
		16'b0000101100101111: color_data = 12'b001110100111;
		16'b0000101100110000: color_data = 12'b001110100111;
		16'b0000101100110001: color_data = 12'b001110100111;
		16'b0000101100110010: color_data = 12'b001110100111;
		16'b0000101100110011: color_data = 12'b001110100111;
		16'b0000101100110100: color_data = 12'b001110100111;
		16'b0000101100110101: color_data = 12'b001110100111;
		16'b0000101100110110: color_data = 12'b001110100111;
		16'b0000101100110111: color_data = 12'b001110100111;
		16'b0000101100111000: color_data = 12'b001110100111;
		16'b0000101100111001: color_data = 12'b001110100111;
		16'b0000101100111010: color_data = 12'b001110100111;
		16'b0000101100111011: color_data = 12'b001110100111;
		16'b0000101100111100: color_data = 12'b001110100111;
		16'b0000101100111101: color_data = 12'b001110100111;
		16'b0000101100111110: color_data = 12'b001110100111;
		16'b0000101100111111: color_data = 12'b001110100111;
		16'b0000101101000000: color_data = 12'b001110100111;
		16'b0000101101000001: color_data = 12'b001110100111;
		16'b0000101101000010: color_data = 12'b001110100111;
		16'b0000101101000011: color_data = 12'b001110100111;
		16'b0000101101000100: color_data = 12'b001110100111;
		16'b0000101101100100: color_data = 12'b001110100111;
		16'b0000101101100101: color_data = 12'b001110100111;
		16'b0000101101100110: color_data = 12'b001110100111;
		16'b0000101101100111: color_data = 12'b001110100111;
		16'b0000101101101000: color_data = 12'b001110100111;
		16'b0000101101101001: color_data = 12'b001110100111;
		16'b0000101101101010: color_data = 12'b001110100111;
		16'b0000101101101011: color_data = 12'b001110100111;
		16'b0000101101101100: color_data = 12'b001110100111;
		16'b0000101101101101: color_data = 12'b001110100111;
		16'b0000101101101110: color_data = 12'b001110100111;
		16'b0000101101101111: color_data = 12'b001110100111;
		16'b0000101101110000: color_data = 12'b001110100111;
		16'b0000101101110001: color_data = 12'b001110100111;
		16'b0000101101110010: color_data = 12'b001110100111;
		16'b0000101101110011: color_data = 12'b001110100111;
		16'b0000101101110100: color_data = 12'b001110100111;
		16'b0000101101110101: color_data = 12'b001110100111;
		16'b0000101101110110: color_data = 12'b001110100111;
		16'b0000101101110111: color_data = 12'b001110100111;
		16'b0000101101111000: color_data = 12'b001110100111;
		16'b0000101101111001: color_data = 12'b001110100111;
		16'b0000101101111010: color_data = 12'b001110100111;
		16'b0000101101111011: color_data = 12'b001110100111;
		16'b0000110000001101: color_data = 12'b001110100111;
		16'b0000110000001110: color_data = 12'b001110100111;
		16'b0000110000001111: color_data = 12'b001110100111;
		16'b0000110000010000: color_data = 12'b001110100111;
		16'b0000110000010001: color_data = 12'b001110100111;
		16'b0000110000010010: color_data = 12'b001110100111;
		16'b0000110000010011: color_data = 12'b001110100111;
		16'b0000110000010100: color_data = 12'b001110100111;
		16'b0000110000010101: color_data = 12'b001110100111;
		16'b0000110000010110: color_data = 12'b001110100111;
		16'b0000110000010111: color_data = 12'b001110100111;
		16'b0000110000011000: color_data = 12'b001110100111;
		16'b0000110000011001: color_data = 12'b001110100111;
		16'b0000110000011010: color_data = 12'b001110100111;
		16'b0000110000011011: color_data = 12'b001110100111;
		16'b0000110000011100: color_data = 12'b001110100111;
		16'b0000110000011101: color_data = 12'b001110100111;
		16'b0000110000011110: color_data = 12'b001110100111;
		16'b0000110000011111: color_data = 12'b001110100111;
		16'b0000110000100000: color_data = 12'b001110100111;
		16'b0000110000100001: color_data = 12'b001110100111;
		16'b0000110000100010: color_data = 12'b001110100111;
		16'b0000110000100011: color_data = 12'b001110100111;
		16'b0000110000100100: color_data = 12'b001110100111;
		16'b0000110000101011: color_data = 12'b001110100111;
		16'b0000110000101100: color_data = 12'b001110100111;
		16'b0000110000101101: color_data = 12'b001110100111;
		16'b0000110000101110: color_data = 12'b001110100111;
		16'b0000110000101111: color_data = 12'b001110100111;
		16'b0000110000110000: color_data = 12'b001110100111;
		16'b0000110000110001: color_data = 12'b001110100111;
		16'b0000110000110010: color_data = 12'b001110100111;
		16'b0000110000110011: color_data = 12'b001110100111;
		16'b0000110000110100: color_data = 12'b001110100111;
		16'b0000110000110101: color_data = 12'b001110100111;
		16'b0000110000110110: color_data = 12'b001110100111;
		16'b0000110000110111: color_data = 12'b001110100111;
		16'b0000110001000100: color_data = 12'b001110100111;
		16'b0000110001000101: color_data = 12'b001110100111;
		16'b0000110001000110: color_data = 12'b001110100111;
		16'b0000110001000111: color_data = 12'b001110100111;
		16'b0000110001001000: color_data = 12'b001110100111;
		16'b0000110001001001: color_data = 12'b001110100111;
		16'b0000110001001010: color_data = 12'b001110100111;
		16'b0000110001001011: color_data = 12'b001110100111;
		16'b0000110001001100: color_data = 12'b001110100111;
		16'b0000110001001101: color_data = 12'b001110100111;
		16'b0000110001001110: color_data = 12'b001110100111;
		16'b0000110001001111: color_data = 12'b001110100111;
		16'b0000110001010110: color_data = 12'b001110100111;
		16'b0000110001010111: color_data = 12'b001110100111;
		16'b0000110001011000: color_data = 12'b001110100111;
		16'b0000110001011001: color_data = 12'b001110100111;
		16'b0000110001011010: color_data = 12'b001110100111;
		16'b0000110001011011: color_data = 12'b001110100111;
		16'b0000110001011100: color_data = 12'b001110100111;
		16'b0000110001011101: color_data = 12'b001110100111;
		16'b0000110001011110: color_data = 12'b001110100111;
		16'b0000110001011111: color_data = 12'b001110100111;
		16'b0000110001100000: color_data = 12'b001110100111;
		16'b0000110001100001: color_data = 12'b001110100111;
		16'b0000110001100010: color_data = 12'b001110100111;
		16'b0000110001100011: color_data = 12'b001110100111;
		16'b0000110001100100: color_data = 12'b001110100111;
		16'b0000110001100101: color_data = 12'b001110100111;
		16'b0000110001100110: color_data = 12'b001110100111;
		16'b0000110001100111: color_data = 12'b001110100111;
		16'b0000110001101000: color_data = 12'b001110100111;
		16'b0000110001101001: color_data = 12'b001110100111;
		16'b0000110001101010: color_data = 12'b001110100111;
		16'b0000110001101011: color_data = 12'b001110100111;
		16'b0000110001101100: color_data = 12'b001110100111;
		16'b0000110001101101: color_data = 12'b001110100111;
		16'b0000110001101110: color_data = 12'b001110100111;
		16'b0000110001110101: color_data = 12'b001110100111;
		16'b0000110001110110: color_data = 12'b001110100111;
		16'b0000110001110111: color_data = 12'b001110100111;
		16'b0000110001111000: color_data = 12'b001110100111;
		16'b0000110001111001: color_data = 12'b001110100111;
		16'b0000110001111010: color_data = 12'b001110100111;
		16'b0000110001111011: color_data = 12'b001110100111;
		16'b0000110001111100: color_data = 12'b001110100111;
		16'b0000110001111101: color_data = 12'b001110100111;
		16'b0000110001111110: color_data = 12'b001110100111;
		16'b0000110001111111: color_data = 12'b001110100111;
		16'b0000110010000000: color_data = 12'b001110100111;
		16'b0000110010000001: color_data = 12'b001110100111;
		16'b0000110010000010: color_data = 12'b001110100111;
		16'b0000110010000011: color_data = 12'b001110100111;
		16'b0000110010000100: color_data = 12'b001110100111;
		16'b0000110010000101: color_data = 12'b001110100111;
		16'b0000110010000110: color_data = 12'b001110100111;
		16'b0000110010000111: color_data = 12'b001110100111;
		16'b0000110010001000: color_data = 12'b001110100111;
		16'b0000110010001001: color_data = 12'b001110100111;
		16'b0000110010001010: color_data = 12'b001110100111;
		16'b0000110010001011: color_data = 12'b001110100111;
		16'b0000110010001100: color_data = 12'b001110100111;
		16'b0000110010101100: color_data = 12'b001110100111;
		16'b0000110010101101: color_data = 12'b001110100111;
		16'b0000110010101110: color_data = 12'b001110100111;
		16'b0000110010101111: color_data = 12'b001110100111;
		16'b0000110010110000: color_data = 12'b001110100111;
		16'b0000110010110001: color_data = 12'b001110100111;
		16'b0000110010110010: color_data = 12'b001110100111;
		16'b0000110010110011: color_data = 12'b001110100111;
		16'b0000110010110100: color_data = 12'b001110100111;
		16'b0000110010110101: color_data = 12'b001110100111;
		16'b0000110010110110: color_data = 12'b001110100111;
		16'b0000110010110111: color_data = 12'b001110100111;
		16'b0000110010111000: color_data = 12'b001110100111;
		16'b0000110010111001: color_data = 12'b001110100111;
		16'b0000110010111010: color_data = 12'b001110100111;
		16'b0000110010111011: color_data = 12'b001110100111;
		16'b0000110010111100: color_data = 12'b001110100111;
		16'b0000110010111101: color_data = 12'b001110100111;
		16'b0000110010111110: color_data = 12'b001110100111;
		16'b0000110010111111: color_data = 12'b001110100111;
		16'b0000110011000000: color_data = 12'b001110100111;
		16'b0000110011000001: color_data = 12'b001110100111;
		16'b0000110011000010: color_data = 12'b001110100111;
		16'b0000110011000011: color_data = 12'b001110100111;
		16'b0000110011000100: color_data = 12'b001110100111;
		16'b0000110011001011: color_data = 12'b001110100111;
		16'b0000110011001100: color_data = 12'b001110100111;
		16'b0000110011001101: color_data = 12'b001110100111;
		16'b0000110011001110: color_data = 12'b001110100111;
		16'b0000110011001111: color_data = 12'b001110100111;
		16'b0000110011010000: color_data = 12'b001110100111;
		16'b0000110011010001: color_data = 12'b001110100111;
		16'b0000110011010010: color_data = 12'b001110100111;
		16'b0000110011010011: color_data = 12'b001110100111;
		16'b0000110011010100: color_data = 12'b001110100111;
		16'b0000110011010101: color_data = 12'b001110100111;
		16'b0000110011010110: color_data = 12'b001110100111;
		16'b0000110011010111: color_data = 12'b001110100111;
		16'b0000110011011000: color_data = 12'b001110100111;
		16'b0000110011011001: color_data = 12'b001110100111;
		16'b0000110011011010: color_data = 12'b001110100111;
		16'b0000110011011011: color_data = 12'b001110100111;
		16'b0000110011011100: color_data = 12'b001110100111;
		16'b0000110011011101: color_data = 12'b001110100111;
		16'b0000110011011110: color_data = 12'b001110100111;
		16'b0000110011011111: color_data = 12'b001110100111;
		16'b0000110011100000: color_data = 12'b001110100111;
		16'b0000110011100001: color_data = 12'b001110100111;
		16'b0000110011100010: color_data = 12'b001110100111;
		16'b0000110011100011: color_data = 12'b001110100111;
		16'b0000110011100100: color_data = 12'b001110100111;
		16'b0000110011100101: color_data = 12'b001110100111;
		16'b0000110011100110: color_data = 12'b001110100111;
		16'b0000110011100111: color_data = 12'b001110100111;
		16'b0000110011101000: color_data = 12'b001110100111;
		16'b0000110011101001: color_data = 12'b001110100111;
		16'b0000110011101010: color_data = 12'b001110100111;
		16'b0000110011101011: color_data = 12'b001110100111;
		16'b0000110011101100: color_data = 12'b001110100111;
		16'b0000110011101101: color_data = 12'b001110100111;
		16'b0000110011101110: color_data = 12'b001110100111;
		16'b0000110011101111: color_data = 12'b001110100111;
		16'b0000110011111100: color_data = 12'b001110100111;
		16'b0000110011111101: color_data = 12'b001110100111;
		16'b0000110011111110: color_data = 12'b001110100111;
		16'b0000110011111111: color_data = 12'b001110100111;
		16'b0000110100000000: color_data = 12'b001110100111;
		16'b0000110100000001: color_data = 12'b001110100111;
		16'b0000110100000010: color_data = 12'b001110100111;
		16'b0000110100000011: color_data = 12'b001110100111;
		16'b0000110100000100: color_data = 12'b001110100111;
		16'b0000110100000101: color_data = 12'b001110100111;
		16'b0000110100000110: color_data = 12'b001110100111;
		16'b0000110100000111: color_data = 12'b001110100111;
		16'b0000110100001000: color_data = 12'b001110100111;
		16'b0000110100001001: color_data = 12'b001110100111;
		16'b0000110100001010: color_data = 12'b001110100111;
		16'b0000110100001011: color_data = 12'b001110100111;
		16'b0000110100001100: color_data = 12'b001110100111;
		16'b0000110100001101: color_data = 12'b001110100111;
		16'b0000110100001110: color_data = 12'b001110100111;
		16'b0000110100001111: color_data = 12'b001110100111;
		16'b0000110100010000: color_data = 12'b001110100111;
		16'b0000110100010001: color_data = 12'b001110100111;
		16'b0000110100010010: color_data = 12'b001110100111;
		16'b0000110100010011: color_data = 12'b001110100111;
		16'b0000110100010100: color_data = 12'b001110100111;
		16'b0000110100010101: color_data = 12'b001110100111;
		16'b0000110100010110: color_data = 12'b001110100111;
		16'b0000110100010111: color_data = 12'b001110100111;
		16'b0000110100011000: color_data = 12'b001110100111;
		16'b0000110100011001: color_data = 12'b001110100111;
		16'b0000110100011010: color_data = 12'b001110100111;
		16'b0000110100011011: color_data = 12'b001110100111;
		16'b0000110100011100: color_data = 12'b001110100111;
		16'b0000110100011101: color_data = 12'b001110100111;
		16'b0000110100011110: color_data = 12'b001110100111;
		16'b0000110100011111: color_data = 12'b001110100111;
		16'b0000110100100000: color_data = 12'b001110100111;
		16'b0000110100101101: color_data = 12'b001110100111;
		16'b0000110100101110: color_data = 12'b001110100111;
		16'b0000110100101111: color_data = 12'b001110100111;
		16'b0000110100110000: color_data = 12'b001110100111;
		16'b0000110100110001: color_data = 12'b001110100111;
		16'b0000110100110010: color_data = 12'b001110100111;
		16'b0000110100110011: color_data = 12'b001110100111;
		16'b0000110100110100: color_data = 12'b001110100111;
		16'b0000110100110101: color_data = 12'b001110100111;
		16'b0000110100110110: color_data = 12'b001110100111;
		16'b0000110100110111: color_data = 12'b001110100111;
		16'b0000110100111000: color_data = 12'b001110100111;
		16'b0000110100111001: color_data = 12'b001110100111;
		16'b0000110100111010: color_data = 12'b001110100111;
		16'b0000110100111011: color_data = 12'b001110100111;
		16'b0000110100111100: color_data = 12'b001110100111;
		16'b0000110100111101: color_data = 12'b001110100111;
		16'b0000110100111110: color_data = 12'b001110100111;
		16'b0000110100111111: color_data = 12'b001110100111;
		16'b0000110101000000: color_data = 12'b001110100111;
		16'b0000110101000001: color_data = 12'b001110100111;
		16'b0000110101000010: color_data = 12'b001110100111;
		16'b0000110101000011: color_data = 12'b001110100111;
		16'b0000110101000100: color_data = 12'b001110100111;
		16'b0000110101100100: color_data = 12'b001110100111;
		16'b0000110101100101: color_data = 12'b001110100111;
		16'b0000110101100110: color_data = 12'b001110100111;
		16'b0000110101100111: color_data = 12'b001110100111;
		16'b0000110101101000: color_data = 12'b001110100111;
		16'b0000110101101001: color_data = 12'b001110100111;
		16'b0000110101101010: color_data = 12'b001110100111;
		16'b0000110101101011: color_data = 12'b001110100111;
		16'b0000110101101100: color_data = 12'b001110100111;
		16'b0000110101101101: color_data = 12'b001110100111;
		16'b0000110101101110: color_data = 12'b001110100111;
		16'b0000110101101111: color_data = 12'b001110100111;
		16'b0000110101110000: color_data = 12'b001110100111;
		16'b0000110101110001: color_data = 12'b001110100111;
		16'b0000110101110010: color_data = 12'b001110100111;
		16'b0000110101110011: color_data = 12'b001110100111;
		16'b0000110101110100: color_data = 12'b001110100111;
		16'b0000110101110101: color_data = 12'b001110100111;
		16'b0000110101110110: color_data = 12'b001110100111;
		16'b0000110101110111: color_data = 12'b001110100111;
		16'b0000110101111000: color_data = 12'b001110100111;
		16'b0000110101111001: color_data = 12'b001110100111;
		16'b0000110101111010: color_data = 12'b001110100111;
		16'b0000110101111011: color_data = 12'b001110100111;
		16'b0000111000001101: color_data = 12'b001110100111;
		16'b0000111000001110: color_data = 12'b001110100111;
		16'b0000111000001111: color_data = 12'b001110100111;
		16'b0000111000010000: color_data = 12'b001110100111;
		16'b0000111000010001: color_data = 12'b001110100111;
		16'b0000111000010010: color_data = 12'b001110100111;
		16'b0000111000010011: color_data = 12'b001110100111;
		16'b0000111000010100: color_data = 12'b001110100111;
		16'b0000111000010101: color_data = 12'b001110100111;
		16'b0000111000010110: color_data = 12'b001110100111;
		16'b0000111000010111: color_data = 12'b001110100111;
		16'b0000111000011000: color_data = 12'b001110100111;
		16'b0000111000011001: color_data = 12'b001110100111;
		16'b0000111000011010: color_data = 12'b001110100111;
		16'b0000111000011011: color_data = 12'b001110100111;
		16'b0000111000011100: color_data = 12'b001110100111;
		16'b0000111000011101: color_data = 12'b001110100111;
		16'b0000111000011110: color_data = 12'b001110100111;
		16'b0000111000011111: color_data = 12'b001110100111;
		16'b0000111000100000: color_data = 12'b001110100111;
		16'b0000111000100001: color_data = 12'b001110100111;
		16'b0000111000100010: color_data = 12'b001110100111;
		16'b0000111000100011: color_data = 12'b001110100111;
		16'b0000111000100100: color_data = 12'b001110100111;
		16'b0000111000101011: color_data = 12'b001110100111;
		16'b0000111000101100: color_data = 12'b001110100111;
		16'b0000111000101101: color_data = 12'b001110100111;
		16'b0000111000101110: color_data = 12'b001110100111;
		16'b0000111000101111: color_data = 12'b001110100111;
		16'b0000111000110000: color_data = 12'b001110100111;
		16'b0000111000110001: color_data = 12'b001110100111;
		16'b0000111000110010: color_data = 12'b001110100111;
		16'b0000111000110011: color_data = 12'b001110100111;
		16'b0000111000110100: color_data = 12'b001110100111;
		16'b0000111000110101: color_data = 12'b001110100111;
		16'b0000111000110110: color_data = 12'b001110100111;
		16'b0000111000110111: color_data = 12'b001110100111;
		16'b0000111001000100: color_data = 12'b001110100111;
		16'b0000111001000101: color_data = 12'b001110100111;
		16'b0000111001000110: color_data = 12'b001110100111;
		16'b0000111001000111: color_data = 12'b001110100111;
		16'b0000111001001000: color_data = 12'b001110100111;
		16'b0000111001001001: color_data = 12'b001110100111;
		16'b0000111001001010: color_data = 12'b001110100111;
		16'b0000111001001011: color_data = 12'b001110100111;
		16'b0000111001001100: color_data = 12'b001110100111;
		16'b0000111001001101: color_data = 12'b001110100111;
		16'b0000111001001110: color_data = 12'b001110100111;
		16'b0000111001001111: color_data = 12'b001110100111;
		16'b0000111001010110: color_data = 12'b001110100111;
		16'b0000111001010111: color_data = 12'b001110100111;
		16'b0000111001011000: color_data = 12'b001110100111;
		16'b0000111001011001: color_data = 12'b001110100111;
		16'b0000111001011010: color_data = 12'b001110100111;
		16'b0000111001011011: color_data = 12'b001110100111;
		16'b0000111001011100: color_data = 12'b001110100111;
		16'b0000111001011101: color_data = 12'b001110100111;
		16'b0000111001011110: color_data = 12'b001110100111;
		16'b0000111001011111: color_data = 12'b001110100111;
		16'b0000111001100000: color_data = 12'b001110100111;
		16'b0000111001100001: color_data = 12'b001110100111;
		16'b0000111001100010: color_data = 12'b001110100111;
		16'b0000111001100011: color_data = 12'b001110100111;
		16'b0000111001100100: color_data = 12'b001110100111;
		16'b0000111001100101: color_data = 12'b001110100111;
		16'b0000111001100110: color_data = 12'b001110100111;
		16'b0000111001100111: color_data = 12'b001110100111;
		16'b0000111001101000: color_data = 12'b001110100111;
		16'b0000111001101001: color_data = 12'b001110100111;
		16'b0000111001101010: color_data = 12'b001110100111;
		16'b0000111001101011: color_data = 12'b001110100111;
		16'b0000111001101100: color_data = 12'b001110100111;
		16'b0000111001101101: color_data = 12'b001110100111;
		16'b0000111001101110: color_data = 12'b001110100111;
		16'b0000111001110101: color_data = 12'b001110100111;
		16'b0000111001110110: color_data = 12'b001110100111;
		16'b0000111001110111: color_data = 12'b001110100111;
		16'b0000111001111000: color_data = 12'b001110100111;
		16'b0000111001111001: color_data = 12'b001110100111;
		16'b0000111001111010: color_data = 12'b001110100111;
		16'b0000111001111011: color_data = 12'b001110100111;
		16'b0000111001111100: color_data = 12'b001110100111;
		16'b0000111001111101: color_data = 12'b001110100111;
		16'b0000111001111110: color_data = 12'b001110100111;
		16'b0000111001111111: color_data = 12'b001110100111;
		16'b0000111010000000: color_data = 12'b001110100111;
		16'b0000111010000001: color_data = 12'b001110100111;
		16'b0000111010000010: color_data = 12'b001110100111;
		16'b0000111010000011: color_data = 12'b001110100111;
		16'b0000111010000100: color_data = 12'b001110100111;
		16'b0000111010000101: color_data = 12'b001110100111;
		16'b0000111010000110: color_data = 12'b001110100111;
		16'b0000111010000111: color_data = 12'b001110100111;
		16'b0000111010001000: color_data = 12'b001110100111;
		16'b0000111010001001: color_data = 12'b001110100111;
		16'b0000111010001010: color_data = 12'b001110100111;
		16'b0000111010001011: color_data = 12'b001110100111;
		16'b0000111010001100: color_data = 12'b001110100111;
		16'b0000111010101100: color_data = 12'b001110100111;
		16'b0000111010101101: color_data = 12'b001110100111;
		16'b0000111010101110: color_data = 12'b001110100111;
		16'b0000111010101111: color_data = 12'b001110100111;
		16'b0000111010110000: color_data = 12'b001110100111;
		16'b0000111010110001: color_data = 12'b001110100111;
		16'b0000111010110010: color_data = 12'b001110100111;
		16'b0000111010110011: color_data = 12'b001110100111;
		16'b0000111010110100: color_data = 12'b001110100111;
		16'b0000111010110101: color_data = 12'b001110100111;
		16'b0000111010110110: color_data = 12'b001110100111;
		16'b0000111010110111: color_data = 12'b001110100111;
		16'b0000111010111000: color_data = 12'b001110100111;
		16'b0000111010111001: color_data = 12'b001110100111;
		16'b0000111010111010: color_data = 12'b001110100111;
		16'b0000111010111011: color_data = 12'b001110100111;
		16'b0000111010111100: color_data = 12'b001110100111;
		16'b0000111010111101: color_data = 12'b001110100111;
		16'b0000111010111110: color_data = 12'b001110100111;
		16'b0000111010111111: color_data = 12'b001110100111;
		16'b0000111011000000: color_data = 12'b001110100111;
		16'b0000111011000001: color_data = 12'b001110100111;
		16'b0000111011000010: color_data = 12'b001110100111;
		16'b0000111011000011: color_data = 12'b001110100111;
		16'b0000111011000100: color_data = 12'b001110100111;
		16'b0000111011001011: color_data = 12'b001110100111;
		16'b0000111011001100: color_data = 12'b001110100111;
		16'b0000111011001101: color_data = 12'b001110100111;
		16'b0000111011001110: color_data = 12'b001110100111;
		16'b0000111011001111: color_data = 12'b001110100111;
		16'b0000111011010000: color_data = 12'b001110100111;
		16'b0000111011010001: color_data = 12'b001110100111;
		16'b0000111011010010: color_data = 12'b001110100111;
		16'b0000111011010011: color_data = 12'b001110100111;
		16'b0000111011010100: color_data = 12'b001110100111;
		16'b0000111011010101: color_data = 12'b001110100111;
		16'b0000111011010110: color_data = 12'b001110100111;
		16'b0000111011010111: color_data = 12'b001110100111;
		16'b0000111011011000: color_data = 12'b001110100111;
		16'b0000111011011001: color_data = 12'b001110100111;
		16'b0000111011011010: color_data = 12'b001110100111;
		16'b0000111011011011: color_data = 12'b001110100111;
		16'b0000111011011100: color_data = 12'b001110100111;
		16'b0000111011011101: color_data = 12'b001110100111;
		16'b0000111011011110: color_data = 12'b001110100111;
		16'b0000111011011111: color_data = 12'b001110100111;
		16'b0000111011100000: color_data = 12'b001110100111;
		16'b0000111011100001: color_data = 12'b001110100111;
		16'b0000111011100010: color_data = 12'b001110100111;
		16'b0000111011100011: color_data = 12'b001110100111;
		16'b0000111011100100: color_data = 12'b001110100111;
		16'b0000111011100101: color_data = 12'b001110100111;
		16'b0000111011100110: color_data = 12'b001110100111;
		16'b0000111011100111: color_data = 12'b001110100111;
		16'b0000111011101000: color_data = 12'b001110100111;
		16'b0000111011101001: color_data = 12'b001110100111;
		16'b0000111011101010: color_data = 12'b001110100111;
		16'b0000111011101011: color_data = 12'b001110100111;
		16'b0000111011101100: color_data = 12'b001110100111;
		16'b0000111011101101: color_data = 12'b001110100111;
		16'b0000111011101110: color_data = 12'b001110100111;
		16'b0000111011101111: color_data = 12'b001110100111;
		16'b0000111011111100: color_data = 12'b001110100111;
		16'b0000111011111101: color_data = 12'b001110100111;
		16'b0000111011111110: color_data = 12'b001110100111;
		16'b0000111011111111: color_data = 12'b001110100111;
		16'b0000111100000000: color_data = 12'b001110100111;
		16'b0000111100000001: color_data = 12'b001110100111;
		16'b0000111100000010: color_data = 12'b001110100111;
		16'b0000111100000011: color_data = 12'b001110100111;
		16'b0000111100000100: color_data = 12'b001110100111;
		16'b0000111100000101: color_data = 12'b001110100111;
		16'b0000111100000110: color_data = 12'b001110100111;
		16'b0000111100000111: color_data = 12'b001110100111;
		16'b0000111100001000: color_data = 12'b001110100111;
		16'b0000111100001001: color_data = 12'b001110100111;
		16'b0000111100001010: color_data = 12'b001110100111;
		16'b0000111100001011: color_data = 12'b001110100111;
		16'b0000111100001100: color_data = 12'b001110100111;
		16'b0000111100001101: color_data = 12'b001110100111;
		16'b0000111100001110: color_data = 12'b001110100111;
		16'b0000111100001111: color_data = 12'b001110100111;
		16'b0000111100010000: color_data = 12'b001110100111;
		16'b0000111100010001: color_data = 12'b001110100111;
		16'b0000111100010010: color_data = 12'b001110100111;
		16'b0000111100010011: color_data = 12'b001110100111;
		16'b0000111100010100: color_data = 12'b001110100111;
		16'b0000111100010101: color_data = 12'b001110100111;
		16'b0000111100010110: color_data = 12'b001110100111;
		16'b0000111100010111: color_data = 12'b001110100111;
		16'b0000111100011000: color_data = 12'b001110100111;
		16'b0000111100011001: color_data = 12'b001110100111;
		16'b0000111100011010: color_data = 12'b001110100111;
		16'b0000111100011011: color_data = 12'b001110100111;
		16'b0000111100011100: color_data = 12'b001110100111;
		16'b0000111100011101: color_data = 12'b001110100111;
		16'b0000111100011110: color_data = 12'b001110100111;
		16'b0000111100011111: color_data = 12'b001110100111;
		16'b0000111100100000: color_data = 12'b001110100111;
		16'b0000111100101101: color_data = 12'b001110100111;
		16'b0000111100101110: color_data = 12'b001110100111;
		16'b0000111100101111: color_data = 12'b001110100111;
		16'b0000111100110000: color_data = 12'b001110100111;
		16'b0000111100110001: color_data = 12'b001110100111;
		16'b0000111100110010: color_data = 12'b001110100111;
		16'b0000111100110011: color_data = 12'b001110100111;
		16'b0000111100110100: color_data = 12'b001110100111;
		16'b0000111100110101: color_data = 12'b001110100111;
		16'b0000111100110110: color_data = 12'b001110100111;
		16'b0000111100110111: color_data = 12'b001110100111;
		16'b0000111100111000: color_data = 12'b001110100111;
		16'b0000111100111001: color_data = 12'b001110100111;
		16'b0000111100111010: color_data = 12'b001110100111;
		16'b0000111100111011: color_data = 12'b001110100111;
		16'b0000111100111100: color_data = 12'b001110100111;
		16'b0000111100111101: color_data = 12'b001110100111;
		16'b0000111100111110: color_data = 12'b001110100111;
		16'b0000111100111111: color_data = 12'b001110100111;
		16'b0000111101000000: color_data = 12'b001110100111;
		16'b0000111101000001: color_data = 12'b001110100111;
		16'b0000111101000010: color_data = 12'b001110100111;
		16'b0000111101000011: color_data = 12'b001110100111;
		16'b0000111101000100: color_data = 12'b001110100111;
		16'b0000111101100100: color_data = 12'b001110100111;
		16'b0000111101100101: color_data = 12'b001110100111;
		16'b0000111101100110: color_data = 12'b001110100111;
		16'b0000111101100111: color_data = 12'b001110100111;
		16'b0000111101101000: color_data = 12'b001110100111;
		16'b0000111101101001: color_data = 12'b001110100111;
		16'b0000111101101010: color_data = 12'b001110100111;
		16'b0000111101101011: color_data = 12'b001110100111;
		16'b0000111101101100: color_data = 12'b001110100111;
		16'b0000111101101101: color_data = 12'b001110100111;
		16'b0000111101101110: color_data = 12'b001110100111;
		16'b0000111101101111: color_data = 12'b001110100111;
		16'b0000111101110000: color_data = 12'b001110100111;
		16'b0000111101110001: color_data = 12'b001110100111;
		16'b0000111101110010: color_data = 12'b001110100111;
		16'b0000111101110011: color_data = 12'b001110100111;
		16'b0000111101110100: color_data = 12'b001110100111;
		16'b0000111101110101: color_data = 12'b001110100111;
		16'b0000111101110110: color_data = 12'b001110100111;
		16'b0000111101110111: color_data = 12'b001110100111;
		16'b0000111101111000: color_data = 12'b001110100111;
		16'b0000111101111001: color_data = 12'b001110100111;
		16'b0000111101111010: color_data = 12'b001110100111;
		16'b0000111101111011: color_data = 12'b001110100111;
		16'b0001000000001101: color_data = 12'b001110100111;
		16'b0001000000001110: color_data = 12'b001110100111;
		16'b0001000000001111: color_data = 12'b001110100111;
		16'b0001000000010000: color_data = 12'b001110100111;
		16'b0001000000010001: color_data = 12'b001110100111;
		16'b0001000000010010: color_data = 12'b001110100111;
		16'b0001000000010011: color_data = 12'b001110100111;
		16'b0001000000010100: color_data = 12'b001110100111;
		16'b0001000000010101: color_data = 12'b001110100111;
		16'b0001000000010110: color_data = 12'b001110100111;
		16'b0001000000010111: color_data = 12'b001110100111;
		16'b0001000000011000: color_data = 12'b001110100111;
		16'b0001000000011001: color_data = 12'b001110100111;
		16'b0001000000011010: color_data = 12'b001110100111;
		16'b0001000000011011: color_data = 12'b001110100111;
		16'b0001000000011100: color_data = 12'b001110100111;
		16'b0001000000011101: color_data = 12'b001110100111;
		16'b0001000000011110: color_data = 12'b001110100111;
		16'b0001000000011111: color_data = 12'b001110100111;
		16'b0001000000100000: color_data = 12'b001110100111;
		16'b0001000000100001: color_data = 12'b001110100111;
		16'b0001000000100010: color_data = 12'b001110100111;
		16'b0001000000100011: color_data = 12'b001110100111;
		16'b0001000000100100: color_data = 12'b001110100111;
		16'b0001000000101011: color_data = 12'b001110100111;
		16'b0001000000101100: color_data = 12'b001110100111;
		16'b0001000000101101: color_data = 12'b001110100111;
		16'b0001000000101110: color_data = 12'b001110100111;
		16'b0001000000101111: color_data = 12'b001110100111;
		16'b0001000000110000: color_data = 12'b001110100111;
		16'b0001000000110001: color_data = 12'b001110100111;
		16'b0001000000110010: color_data = 12'b001110100111;
		16'b0001000000110011: color_data = 12'b001110100111;
		16'b0001000000110100: color_data = 12'b001110100111;
		16'b0001000000110101: color_data = 12'b001110100111;
		16'b0001000000110110: color_data = 12'b001110100111;
		16'b0001000000110111: color_data = 12'b001110100111;
		16'b0001000001000100: color_data = 12'b001110100111;
		16'b0001000001000101: color_data = 12'b001110100111;
		16'b0001000001000110: color_data = 12'b001110100111;
		16'b0001000001000111: color_data = 12'b001110100111;
		16'b0001000001001000: color_data = 12'b001110100111;
		16'b0001000001001001: color_data = 12'b001110100111;
		16'b0001000001001010: color_data = 12'b001110100111;
		16'b0001000001001011: color_data = 12'b001110100111;
		16'b0001000001001100: color_data = 12'b001110100111;
		16'b0001000001001101: color_data = 12'b001110100111;
		16'b0001000001001110: color_data = 12'b001110100111;
		16'b0001000001001111: color_data = 12'b001110100111;
		16'b0001000001010110: color_data = 12'b001110100111;
		16'b0001000001010111: color_data = 12'b001110100111;
		16'b0001000001011000: color_data = 12'b001110100111;
		16'b0001000001011001: color_data = 12'b001110100111;
		16'b0001000001011010: color_data = 12'b001110100111;
		16'b0001000001011011: color_data = 12'b001110100111;
		16'b0001000001011100: color_data = 12'b001110100111;
		16'b0001000001011101: color_data = 12'b001110100111;
		16'b0001000001011110: color_data = 12'b001110100111;
		16'b0001000001011111: color_data = 12'b001110100111;
		16'b0001000001100000: color_data = 12'b001110100111;
		16'b0001000001100001: color_data = 12'b001110100111;
		16'b0001000001100010: color_data = 12'b001110100111;
		16'b0001000001100011: color_data = 12'b001110100111;
		16'b0001000001100100: color_data = 12'b001110100111;
		16'b0001000001100101: color_data = 12'b001110100111;
		16'b0001000001100110: color_data = 12'b001110100111;
		16'b0001000001100111: color_data = 12'b001110100111;
		16'b0001000001101000: color_data = 12'b001110100111;
		16'b0001000001101001: color_data = 12'b001110100111;
		16'b0001000001101010: color_data = 12'b001110100111;
		16'b0001000001101011: color_data = 12'b001110100111;
		16'b0001000001101100: color_data = 12'b001110100111;
		16'b0001000001101101: color_data = 12'b001110100111;
		16'b0001000001101110: color_data = 12'b001110100111;
		16'b0001000001110101: color_data = 12'b001110100111;
		16'b0001000001110110: color_data = 12'b001110100111;
		16'b0001000001110111: color_data = 12'b001110100111;
		16'b0001000001111000: color_data = 12'b001110100111;
		16'b0001000001111001: color_data = 12'b001110100111;
		16'b0001000001111010: color_data = 12'b001110100111;
		16'b0001000001111011: color_data = 12'b001110100111;
		16'b0001000001111100: color_data = 12'b001110100111;
		16'b0001000001111101: color_data = 12'b001110100111;
		16'b0001000001111110: color_data = 12'b001110100111;
		16'b0001000001111111: color_data = 12'b001110100111;
		16'b0001000010000000: color_data = 12'b001110100111;
		16'b0001000010000001: color_data = 12'b001110100111;
		16'b0001000010000010: color_data = 12'b001110100111;
		16'b0001000010000011: color_data = 12'b001110100111;
		16'b0001000010000100: color_data = 12'b001110100111;
		16'b0001000010000101: color_data = 12'b001110100111;
		16'b0001000010000110: color_data = 12'b001110100111;
		16'b0001000010000111: color_data = 12'b001110100111;
		16'b0001000010001000: color_data = 12'b001110100111;
		16'b0001000010001001: color_data = 12'b001110100111;
		16'b0001000010001010: color_data = 12'b001110100111;
		16'b0001000010001011: color_data = 12'b001110100111;
		16'b0001000010001100: color_data = 12'b001110100111;
		16'b0001000010101100: color_data = 12'b001110100111;
		16'b0001000010101101: color_data = 12'b001110100111;
		16'b0001000010101110: color_data = 12'b001110100111;
		16'b0001000010101111: color_data = 12'b001110100111;
		16'b0001000010110000: color_data = 12'b001110100111;
		16'b0001000010110001: color_data = 12'b001110100111;
		16'b0001000010110010: color_data = 12'b001110100111;
		16'b0001000010110011: color_data = 12'b001110100111;
		16'b0001000010110100: color_data = 12'b001110100111;
		16'b0001000010110101: color_data = 12'b001110100111;
		16'b0001000010110110: color_data = 12'b001110100111;
		16'b0001000010110111: color_data = 12'b001110100111;
		16'b0001000010111000: color_data = 12'b001110100111;
		16'b0001000010111001: color_data = 12'b001110100111;
		16'b0001000010111010: color_data = 12'b001110100111;
		16'b0001000010111011: color_data = 12'b001110100111;
		16'b0001000010111100: color_data = 12'b001110100111;
		16'b0001000010111101: color_data = 12'b001110100111;
		16'b0001000010111110: color_data = 12'b001110100111;
		16'b0001000010111111: color_data = 12'b001110100111;
		16'b0001000011000000: color_data = 12'b001110100111;
		16'b0001000011000001: color_data = 12'b001110100111;
		16'b0001000011000010: color_data = 12'b001110100111;
		16'b0001000011000011: color_data = 12'b001110100111;
		16'b0001000011000100: color_data = 12'b001110100111;
		16'b0001000011001011: color_data = 12'b001110100111;
		16'b0001000011001100: color_data = 12'b001110100111;
		16'b0001000011001101: color_data = 12'b001110100111;
		16'b0001000011001110: color_data = 12'b001110100111;
		16'b0001000011001111: color_data = 12'b001110100111;
		16'b0001000011010000: color_data = 12'b001110100111;
		16'b0001000011010001: color_data = 12'b001110100111;
		16'b0001000011010010: color_data = 12'b001110100111;
		16'b0001000011010011: color_data = 12'b001110100111;
		16'b0001000011010100: color_data = 12'b001110100111;
		16'b0001000011010101: color_data = 12'b001110100111;
		16'b0001000011010110: color_data = 12'b001110100111;
		16'b0001000011010111: color_data = 12'b001110100111;
		16'b0001000011011000: color_data = 12'b001110100111;
		16'b0001000011011001: color_data = 12'b001110100111;
		16'b0001000011011010: color_data = 12'b001110100111;
		16'b0001000011011011: color_data = 12'b001110100111;
		16'b0001000011011100: color_data = 12'b001110100111;
		16'b0001000011011101: color_data = 12'b001110100111;
		16'b0001000011011110: color_data = 12'b001110100111;
		16'b0001000011011111: color_data = 12'b001110100111;
		16'b0001000011100000: color_data = 12'b001110100111;
		16'b0001000011100001: color_data = 12'b001110100111;
		16'b0001000011100010: color_data = 12'b001110100111;
		16'b0001000011100011: color_data = 12'b001110100111;
		16'b0001000011100100: color_data = 12'b001110100111;
		16'b0001000011100101: color_data = 12'b001110100111;
		16'b0001000011100110: color_data = 12'b001110100111;
		16'b0001000011100111: color_data = 12'b001110100111;
		16'b0001000011101000: color_data = 12'b001110100111;
		16'b0001000011101001: color_data = 12'b001110100111;
		16'b0001000011101010: color_data = 12'b001110100111;
		16'b0001000011101011: color_data = 12'b001110100111;
		16'b0001000011101100: color_data = 12'b001110100111;
		16'b0001000011101101: color_data = 12'b001110100111;
		16'b0001000011101110: color_data = 12'b001110100111;
		16'b0001000011101111: color_data = 12'b001110100111;
		16'b0001000011111100: color_data = 12'b001110100111;
		16'b0001000011111101: color_data = 12'b001110100111;
		16'b0001000011111110: color_data = 12'b001110100111;
		16'b0001000011111111: color_data = 12'b001110100111;
		16'b0001000100000000: color_data = 12'b001110100111;
		16'b0001000100000001: color_data = 12'b001110100111;
		16'b0001000100000010: color_data = 12'b001110100111;
		16'b0001000100000011: color_data = 12'b001110100111;
		16'b0001000100000100: color_data = 12'b001110100111;
		16'b0001000100000101: color_data = 12'b001110100111;
		16'b0001000100000110: color_data = 12'b001110100111;
		16'b0001000100000111: color_data = 12'b001110100111;
		16'b0001000100001000: color_data = 12'b001110100111;
		16'b0001000100001001: color_data = 12'b001110100111;
		16'b0001000100001010: color_data = 12'b001110100111;
		16'b0001000100001011: color_data = 12'b001110100111;
		16'b0001000100001100: color_data = 12'b001110100111;
		16'b0001000100001101: color_data = 12'b001110100111;
		16'b0001000100001110: color_data = 12'b001110100111;
		16'b0001000100001111: color_data = 12'b001110100111;
		16'b0001000100010000: color_data = 12'b001110100111;
		16'b0001000100010001: color_data = 12'b001110100111;
		16'b0001000100010010: color_data = 12'b001110100111;
		16'b0001000100010011: color_data = 12'b001110100111;
		16'b0001000100010100: color_data = 12'b001110100111;
		16'b0001000100010101: color_data = 12'b001110100111;
		16'b0001000100010110: color_data = 12'b001110100111;
		16'b0001000100010111: color_data = 12'b001110100111;
		16'b0001000100011000: color_data = 12'b001110100111;
		16'b0001000100011001: color_data = 12'b001110100111;
		16'b0001000100011010: color_data = 12'b001110100111;
		16'b0001000100011011: color_data = 12'b001110100111;
		16'b0001000100011100: color_data = 12'b001110100111;
		16'b0001000100011101: color_data = 12'b001110100111;
		16'b0001000100011110: color_data = 12'b001110100111;
		16'b0001000100011111: color_data = 12'b001110100111;
		16'b0001000100100000: color_data = 12'b001110100111;
		16'b0001000100101101: color_data = 12'b001110100111;
		16'b0001000100101110: color_data = 12'b001110100111;
		16'b0001000100101111: color_data = 12'b001110100111;
		16'b0001000100110000: color_data = 12'b001110100111;
		16'b0001000100110001: color_data = 12'b001110100111;
		16'b0001000100110010: color_data = 12'b001110100111;
		16'b0001000100110011: color_data = 12'b001110100111;
		16'b0001000100110100: color_data = 12'b001110100111;
		16'b0001000100110101: color_data = 12'b001110100111;
		16'b0001000100110110: color_data = 12'b001110100111;
		16'b0001000100110111: color_data = 12'b001110100111;
		16'b0001000100111000: color_data = 12'b001110100111;
		16'b0001000100111001: color_data = 12'b001110100111;
		16'b0001000100111010: color_data = 12'b001110100111;
		16'b0001000100111011: color_data = 12'b001110100111;
		16'b0001000100111100: color_data = 12'b001110100111;
		16'b0001000100111101: color_data = 12'b001110100111;
		16'b0001000100111110: color_data = 12'b001110100111;
		16'b0001000100111111: color_data = 12'b001110100111;
		16'b0001000101000000: color_data = 12'b001110100111;
		16'b0001000101000001: color_data = 12'b001110100111;
		16'b0001000101000010: color_data = 12'b001110100111;
		16'b0001000101000011: color_data = 12'b001110100111;
		16'b0001000101000100: color_data = 12'b001110100111;
		16'b0001000101100100: color_data = 12'b001110100111;
		16'b0001000101100101: color_data = 12'b001110100111;
		16'b0001000101100110: color_data = 12'b001110100111;
		16'b0001000101100111: color_data = 12'b001110100111;
		16'b0001000101101000: color_data = 12'b001110100111;
		16'b0001000101101001: color_data = 12'b001110100111;
		16'b0001000101101010: color_data = 12'b001110100111;
		16'b0001000101101011: color_data = 12'b001110100111;
		16'b0001000101101100: color_data = 12'b001110100111;
		16'b0001000101101101: color_data = 12'b001110100111;
		16'b0001000101101110: color_data = 12'b001110100111;
		16'b0001000101101111: color_data = 12'b001110100111;
		16'b0001000101110000: color_data = 12'b001110100111;
		16'b0001000101110001: color_data = 12'b001110100111;
		16'b0001000101110010: color_data = 12'b001110100111;
		16'b0001000101110011: color_data = 12'b001110100111;
		16'b0001000101110100: color_data = 12'b001110100111;
		16'b0001000101110101: color_data = 12'b001110100111;
		16'b0001000101110110: color_data = 12'b001110100111;
		16'b0001000101110111: color_data = 12'b001110100111;
		16'b0001000101111000: color_data = 12'b001110100111;
		16'b0001000101111001: color_data = 12'b001110100111;
		16'b0001000101111010: color_data = 12'b001110100111;
		16'b0001000101111011: color_data = 12'b001110100111;
		16'b0001001000001101: color_data = 12'b001110100111;
		16'b0001001000001110: color_data = 12'b001110100111;
		16'b0001001000001111: color_data = 12'b001110100111;
		16'b0001001000010000: color_data = 12'b001110100111;
		16'b0001001000010001: color_data = 12'b001110100111;
		16'b0001001000010010: color_data = 12'b001110100111;
		16'b0001001000010011: color_data = 12'b001110100111;
		16'b0001001000010100: color_data = 12'b001110100111;
		16'b0001001000010101: color_data = 12'b001110100111;
		16'b0001001000010110: color_data = 12'b001110100111;
		16'b0001001000010111: color_data = 12'b001110100111;
		16'b0001001000011000: color_data = 12'b001110100111;
		16'b0001001000011001: color_data = 12'b001110100111;
		16'b0001001000011010: color_data = 12'b001110100111;
		16'b0001001000011011: color_data = 12'b001110100111;
		16'b0001001000011100: color_data = 12'b001110100111;
		16'b0001001000011101: color_data = 12'b001110100111;
		16'b0001001000011110: color_data = 12'b001110100111;
		16'b0001001000011111: color_data = 12'b001110100111;
		16'b0001001000100000: color_data = 12'b001110100111;
		16'b0001001000100001: color_data = 12'b001110100111;
		16'b0001001000100010: color_data = 12'b001110100111;
		16'b0001001000100011: color_data = 12'b001110100111;
		16'b0001001000100100: color_data = 12'b001110100111;
		16'b0001001000101011: color_data = 12'b001110100111;
		16'b0001001000101100: color_data = 12'b001110100111;
		16'b0001001000101101: color_data = 12'b001110100111;
		16'b0001001000101110: color_data = 12'b001110100111;
		16'b0001001000101111: color_data = 12'b001110100111;
		16'b0001001000110000: color_data = 12'b001110100111;
		16'b0001001000110001: color_data = 12'b001110100111;
		16'b0001001000110010: color_data = 12'b001110100111;
		16'b0001001000110011: color_data = 12'b001110100111;
		16'b0001001000110100: color_data = 12'b001110100111;
		16'b0001001000110101: color_data = 12'b001110100111;
		16'b0001001000110110: color_data = 12'b001110100111;
		16'b0001001000110111: color_data = 12'b001110100111;
		16'b0001001001000100: color_data = 12'b001110100111;
		16'b0001001001000101: color_data = 12'b001110100111;
		16'b0001001001000110: color_data = 12'b001110100111;
		16'b0001001001000111: color_data = 12'b001110100111;
		16'b0001001001001000: color_data = 12'b001110100111;
		16'b0001001001001001: color_data = 12'b001110100111;
		16'b0001001001001010: color_data = 12'b001110100111;
		16'b0001001001001011: color_data = 12'b001110100111;
		16'b0001001001001100: color_data = 12'b001110100111;
		16'b0001001001001101: color_data = 12'b001110100111;
		16'b0001001001001110: color_data = 12'b001110100111;
		16'b0001001001001111: color_data = 12'b001110100111;
		16'b0001001001010110: color_data = 12'b001110100111;
		16'b0001001001010111: color_data = 12'b001110100111;
		16'b0001001001011000: color_data = 12'b001110100111;
		16'b0001001001011001: color_data = 12'b001110100111;
		16'b0001001001011010: color_data = 12'b001110100111;
		16'b0001001001011011: color_data = 12'b001110100111;
		16'b0001001001011100: color_data = 12'b001110100111;
		16'b0001001001011101: color_data = 12'b001110100111;
		16'b0001001001011110: color_data = 12'b001110100111;
		16'b0001001001011111: color_data = 12'b001110100111;
		16'b0001001001100000: color_data = 12'b001110100111;
		16'b0001001001100001: color_data = 12'b001110100111;
		16'b0001001001100010: color_data = 12'b001110100111;
		16'b0001001001100011: color_data = 12'b001110100111;
		16'b0001001001100100: color_data = 12'b001110100111;
		16'b0001001001100101: color_data = 12'b001110100111;
		16'b0001001001100110: color_data = 12'b001110100111;
		16'b0001001001100111: color_data = 12'b001110100111;
		16'b0001001001101000: color_data = 12'b001110100111;
		16'b0001001001101001: color_data = 12'b001110100111;
		16'b0001001001101010: color_data = 12'b001110100111;
		16'b0001001001101011: color_data = 12'b001110100111;
		16'b0001001001101100: color_data = 12'b001110100111;
		16'b0001001001101101: color_data = 12'b001110100111;
		16'b0001001001101110: color_data = 12'b001110100111;
		16'b0001001001110101: color_data = 12'b001110100111;
		16'b0001001001110110: color_data = 12'b001110100111;
		16'b0001001001110111: color_data = 12'b001110100111;
		16'b0001001001111000: color_data = 12'b001110100111;
		16'b0001001001111001: color_data = 12'b001110100111;
		16'b0001001001111010: color_data = 12'b001110100111;
		16'b0001001001111011: color_data = 12'b001110100111;
		16'b0001001001111100: color_data = 12'b001110100111;
		16'b0001001001111101: color_data = 12'b001110100111;
		16'b0001001001111110: color_data = 12'b001110100111;
		16'b0001001001111111: color_data = 12'b001110100111;
		16'b0001001010000000: color_data = 12'b001110100111;
		16'b0001001010000001: color_data = 12'b001110100111;
		16'b0001001010000010: color_data = 12'b001110100111;
		16'b0001001010000011: color_data = 12'b001110100111;
		16'b0001001010000100: color_data = 12'b001110100111;
		16'b0001001010000101: color_data = 12'b001110100111;
		16'b0001001010000110: color_data = 12'b001110100111;
		16'b0001001010000111: color_data = 12'b001110100111;
		16'b0001001010001000: color_data = 12'b001110100111;
		16'b0001001010001001: color_data = 12'b001110100111;
		16'b0001001010001010: color_data = 12'b001110100111;
		16'b0001001010001011: color_data = 12'b001110100111;
		16'b0001001010001100: color_data = 12'b001110100111;
		16'b0001001010101100: color_data = 12'b001110100111;
		16'b0001001010101101: color_data = 12'b001110100111;
		16'b0001001010101110: color_data = 12'b001110100111;
		16'b0001001010101111: color_data = 12'b001110100111;
		16'b0001001010110000: color_data = 12'b001110100111;
		16'b0001001010110001: color_data = 12'b001110100111;
		16'b0001001010110010: color_data = 12'b001110100111;
		16'b0001001010110011: color_data = 12'b001110100111;
		16'b0001001010110100: color_data = 12'b001110100111;
		16'b0001001010110101: color_data = 12'b001110100111;
		16'b0001001010110110: color_data = 12'b001110100111;
		16'b0001001010110111: color_data = 12'b001110100111;
		16'b0001001010111000: color_data = 12'b001110100111;
		16'b0001001010111001: color_data = 12'b001110100111;
		16'b0001001010111010: color_data = 12'b001110100111;
		16'b0001001010111011: color_data = 12'b001110100111;
		16'b0001001010111100: color_data = 12'b001110100111;
		16'b0001001010111101: color_data = 12'b001110100111;
		16'b0001001010111110: color_data = 12'b001110100111;
		16'b0001001010111111: color_data = 12'b001110100111;
		16'b0001001011000000: color_data = 12'b001110100111;
		16'b0001001011000001: color_data = 12'b001110100111;
		16'b0001001011000010: color_data = 12'b001110100111;
		16'b0001001011000011: color_data = 12'b001110100111;
		16'b0001001011000100: color_data = 12'b001110100111;
		16'b0001001011001011: color_data = 12'b001110100111;
		16'b0001001011001100: color_data = 12'b001110100111;
		16'b0001001011001101: color_data = 12'b001110100111;
		16'b0001001011001110: color_data = 12'b001110100111;
		16'b0001001011001111: color_data = 12'b001110100111;
		16'b0001001011010000: color_data = 12'b001110100111;
		16'b0001001011010001: color_data = 12'b001110100111;
		16'b0001001011010010: color_data = 12'b001110100111;
		16'b0001001011010011: color_data = 12'b001110100111;
		16'b0001001011010100: color_data = 12'b001110100111;
		16'b0001001011010101: color_data = 12'b001110100111;
		16'b0001001011010110: color_data = 12'b001110100111;
		16'b0001001011010111: color_data = 12'b001110100111;
		16'b0001001011011000: color_data = 12'b001110100111;
		16'b0001001011011001: color_data = 12'b001110100111;
		16'b0001001011011010: color_data = 12'b001110100111;
		16'b0001001011011011: color_data = 12'b001110100111;
		16'b0001001011011100: color_data = 12'b001110100111;
		16'b0001001011011101: color_data = 12'b001110100111;
		16'b0001001011011110: color_data = 12'b001110100111;
		16'b0001001011011111: color_data = 12'b001110100111;
		16'b0001001011100000: color_data = 12'b001110100111;
		16'b0001001011100001: color_data = 12'b001110100111;
		16'b0001001011100010: color_data = 12'b001110100111;
		16'b0001001011100011: color_data = 12'b001110100111;
		16'b0001001011100100: color_data = 12'b001110100111;
		16'b0001001011100101: color_data = 12'b001110100111;
		16'b0001001011100110: color_data = 12'b001110100111;
		16'b0001001011100111: color_data = 12'b001110100111;
		16'b0001001011101000: color_data = 12'b001110100111;
		16'b0001001011101001: color_data = 12'b001110100111;
		16'b0001001011101010: color_data = 12'b001110100111;
		16'b0001001011101011: color_data = 12'b001110100111;
		16'b0001001011101100: color_data = 12'b001110100111;
		16'b0001001011101101: color_data = 12'b001110100111;
		16'b0001001011101110: color_data = 12'b001110100111;
		16'b0001001011101111: color_data = 12'b001110100111;
		16'b0001001011111100: color_data = 12'b001110100111;
		16'b0001001011111101: color_data = 12'b001110100111;
		16'b0001001011111110: color_data = 12'b001110100111;
		16'b0001001011111111: color_data = 12'b001110100111;
		16'b0001001100000000: color_data = 12'b001110100111;
		16'b0001001100000001: color_data = 12'b001110100111;
		16'b0001001100000010: color_data = 12'b001110100111;
		16'b0001001100000011: color_data = 12'b001110100111;
		16'b0001001100000100: color_data = 12'b001110100111;
		16'b0001001100000101: color_data = 12'b001110100111;
		16'b0001001100000110: color_data = 12'b001110100111;
		16'b0001001100000111: color_data = 12'b001110100111;
		16'b0001001100001000: color_data = 12'b001110100111;
		16'b0001001100001001: color_data = 12'b001110100111;
		16'b0001001100001010: color_data = 12'b001110100111;
		16'b0001001100001011: color_data = 12'b001110100111;
		16'b0001001100001100: color_data = 12'b001110100111;
		16'b0001001100001101: color_data = 12'b001110100111;
		16'b0001001100001110: color_data = 12'b001110100111;
		16'b0001001100001111: color_data = 12'b001110100111;
		16'b0001001100010000: color_data = 12'b001110100111;
		16'b0001001100010001: color_data = 12'b001110100111;
		16'b0001001100010010: color_data = 12'b001110100111;
		16'b0001001100010011: color_data = 12'b001110100111;
		16'b0001001100010100: color_data = 12'b001110100111;
		16'b0001001100010101: color_data = 12'b001110100111;
		16'b0001001100010110: color_data = 12'b001110100111;
		16'b0001001100010111: color_data = 12'b001110100111;
		16'b0001001100011000: color_data = 12'b001110100111;
		16'b0001001100011001: color_data = 12'b001110100111;
		16'b0001001100011010: color_data = 12'b001110100111;
		16'b0001001100011011: color_data = 12'b001110100111;
		16'b0001001100011100: color_data = 12'b001110100111;
		16'b0001001100011101: color_data = 12'b001110100111;
		16'b0001001100011110: color_data = 12'b001110100111;
		16'b0001001100011111: color_data = 12'b001110100111;
		16'b0001001100100000: color_data = 12'b001110100111;
		16'b0001001100101101: color_data = 12'b001110100111;
		16'b0001001100101110: color_data = 12'b001110100111;
		16'b0001001100101111: color_data = 12'b001110100111;
		16'b0001001100110000: color_data = 12'b001110100111;
		16'b0001001100110001: color_data = 12'b001110100111;
		16'b0001001100110010: color_data = 12'b001110100111;
		16'b0001001100110011: color_data = 12'b001110100111;
		16'b0001001100110100: color_data = 12'b001110100111;
		16'b0001001100110101: color_data = 12'b001110100111;
		16'b0001001100110110: color_data = 12'b001110100111;
		16'b0001001100110111: color_data = 12'b001110100111;
		16'b0001001100111000: color_data = 12'b001110100111;
		16'b0001001100111001: color_data = 12'b001110100111;
		16'b0001001100111010: color_data = 12'b001110100111;
		16'b0001001100111011: color_data = 12'b001110100111;
		16'b0001001100111100: color_data = 12'b001110100111;
		16'b0001001100111101: color_data = 12'b001110100111;
		16'b0001001100111110: color_data = 12'b001110100111;
		16'b0001001100111111: color_data = 12'b001110100111;
		16'b0001001101000000: color_data = 12'b001110100111;
		16'b0001001101000001: color_data = 12'b001110100111;
		16'b0001001101000010: color_data = 12'b001110100111;
		16'b0001001101000011: color_data = 12'b001110100111;
		16'b0001001101000100: color_data = 12'b001110100111;
		16'b0001001101100100: color_data = 12'b001110100111;
		16'b0001001101100101: color_data = 12'b001110100111;
		16'b0001001101100110: color_data = 12'b001110100111;
		16'b0001001101100111: color_data = 12'b001110100111;
		16'b0001001101101000: color_data = 12'b001110100111;
		16'b0001001101101001: color_data = 12'b001110100111;
		16'b0001001101101010: color_data = 12'b001110100111;
		16'b0001001101101011: color_data = 12'b001110100111;
		16'b0001001101101100: color_data = 12'b001110100111;
		16'b0001001101101101: color_data = 12'b001110100111;
		16'b0001001101101110: color_data = 12'b001110100111;
		16'b0001001101101111: color_data = 12'b001110100111;
		16'b0001001101110000: color_data = 12'b001110100111;
		16'b0001001101110001: color_data = 12'b001110100111;
		16'b0001001101110010: color_data = 12'b001110100111;
		16'b0001001101110011: color_data = 12'b001110100111;
		16'b0001001101110100: color_data = 12'b001110100111;
		16'b0001001101110101: color_data = 12'b001110100111;
		16'b0001001101110110: color_data = 12'b001110100111;
		16'b0001001101110111: color_data = 12'b001110100111;
		16'b0001001101111000: color_data = 12'b001110100111;
		16'b0001001101111001: color_data = 12'b001110100111;
		16'b0001001101111010: color_data = 12'b001110100111;
		16'b0001001101111011: color_data = 12'b001110100111;
		16'b0001010000001101: color_data = 12'b001110100111;
		16'b0001010000001110: color_data = 12'b001110100111;
		16'b0001010000001111: color_data = 12'b001110100111;
		16'b0001010000010000: color_data = 12'b001110100111;
		16'b0001010000010001: color_data = 12'b001110100111;
		16'b0001010000010010: color_data = 12'b001110100111;
		16'b0001010000010011: color_data = 12'b001110100111;
		16'b0001010000010100: color_data = 12'b001110100111;
		16'b0001010000010101: color_data = 12'b001110100111;
		16'b0001010000010110: color_data = 12'b001110100111;
		16'b0001010000010111: color_data = 12'b001110100111;
		16'b0001010000011000: color_data = 12'b001110100111;
		16'b0001010000011001: color_data = 12'b001110100111;
		16'b0001010000011010: color_data = 12'b001110100111;
		16'b0001010000011011: color_data = 12'b001110100111;
		16'b0001010000011100: color_data = 12'b001110100111;
		16'b0001010000011101: color_data = 12'b001110100111;
		16'b0001010000011110: color_data = 12'b001110100111;
		16'b0001010000011111: color_data = 12'b001110100111;
		16'b0001010000100000: color_data = 12'b001110100111;
		16'b0001010000100001: color_data = 12'b001110100111;
		16'b0001010000100010: color_data = 12'b001110100111;
		16'b0001010000100011: color_data = 12'b001110100111;
		16'b0001010000100100: color_data = 12'b001110100111;
		16'b0001010000101011: color_data = 12'b001110100111;
		16'b0001010000101100: color_data = 12'b001110100111;
		16'b0001010000101101: color_data = 12'b001110100111;
		16'b0001010000101110: color_data = 12'b001110100111;
		16'b0001010000101111: color_data = 12'b001110100111;
		16'b0001010000110000: color_data = 12'b001110100111;
		16'b0001010000110001: color_data = 12'b001110100111;
		16'b0001010000110010: color_data = 12'b001110100111;
		16'b0001010000110011: color_data = 12'b001110100111;
		16'b0001010000110100: color_data = 12'b001110100111;
		16'b0001010000110101: color_data = 12'b001110100111;
		16'b0001010000110110: color_data = 12'b001110100111;
		16'b0001010000110111: color_data = 12'b001110100111;
		16'b0001010001000100: color_data = 12'b001110100111;
		16'b0001010001000101: color_data = 12'b001110100111;
		16'b0001010001000110: color_data = 12'b001110100111;
		16'b0001010001000111: color_data = 12'b001110100111;
		16'b0001010001001000: color_data = 12'b001110100111;
		16'b0001010001001001: color_data = 12'b001110100111;
		16'b0001010001001010: color_data = 12'b001110100111;
		16'b0001010001001011: color_data = 12'b001110100111;
		16'b0001010001001100: color_data = 12'b001110100111;
		16'b0001010001001101: color_data = 12'b001110100111;
		16'b0001010001001110: color_data = 12'b001110100111;
		16'b0001010001001111: color_data = 12'b001110100111;
		16'b0001010001010110: color_data = 12'b001110100111;
		16'b0001010001010111: color_data = 12'b001110100111;
		16'b0001010001011000: color_data = 12'b001110100111;
		16'b0001010001011001: color_data = 12'b001110100111;
		16'b0001010001011010: color_data = 12'b001110100111;
		16'b0001010001011011: color_data = 12'b001110100111;
		16'b0001010001011100: color_data = 12'b001110100111;
		16'b0001010001011101: color_data = 12'b001110100111;
		16'b0001010001011110: color_data = 12'b001110100111;
		16'b0001010001011111: color_data = 12'b001110100111;
		16'b0001010001100000: color_data = 12'b001110100111;
		16'b0001010001100001: color_data = 12'b001110100111;
		16'b0001010001100010: color_data = 12'b001110100111;
		16'b0001010001100011: color_data = 12'b001110100111;
		16'b0001010001100100: color_data = 12'b001110100111;
		16'b0001010001100101: color_data = 12'b001110100111;
		16'b0001010001100110: color_data = 12'b001110100111;
		16'b0001010001100111: color_data = 12'b001110100111;
		16'b0001010001101000: color_data = 12'b001110100111;
		16'b0001010001101001: color_data = 12'b001110100111;
		16'b0001010001101010: color_data = 12'b001110100111;
		16'b0001010001101011: color_data = 12'b001110100111;
		16'b0001010001101100: color_data = 12'b001110100111;
		16'b0001010001101101: color_data = 12'b001110100111;
		16'b0001010001101110: color_data = 12'b001110100111;
		16'b0001010001110101: color_data = 12'b001110100111;
		16'b0001010001110110: color_data = 12'b001110100111;
		16'b0001010001110111: color_data = 12'b001110100111;
		16'b0001010001111000: color_data = 12'b001110100111;
		16'b0001010001111001: color_data = 12'b001110100111;
		16'b0001010001111010: color_data = 12'b001110100111;
		16'b0001010001111011: color_data = 12'b001110100111;
		16'b0001010001111100: color_data = 12'b001110100111;
		16'b0001010001111101: color_data = 12'b001110100111;
		16'b0001010001111110: color_data = 12'b001110100111;
		16'b0001010001111111: color_data = 12'b001110100111;
		16'b0001010010000000: color_data = 12'b001110100111;
		16'b0001010010000001: color_data = 12'b001110100111;
		16'b0001010010000010: color_data = 12'b001110100111;
		16'b0001010010000011: color_data = 12'b001110100111;
		16'b0001010010000100: color_data = 12'b001110100111;
		16'b0001010010000101: color_data = 12'b001110100111;
		16'b0001010010000110: color_data = 12'b001110100111;
		16'b0001010010000111: color_data = 12'b001110100111;
		16'b0001010010001000: color_data = 12'b001110100111;
		16'b0001010010001001: color_data = 12'b001110100111;
		16'b0001010010001010: color_data = 12'b001110100111;
		16'b0001010010001011: color_data = 12'b001110100111;
		16'b0001010010001100: color_data = 12'b001110100111;
		16'b0001010010101100: color_data = 12'b001110100111;
		16'b0001010010101101: color_data = 12'b001110100111;
		16'b0001010010101110: color_data = 12'b001110100111;
		16'b0001010010101111: color_data = 12'b001110100111;
		16'b0001010010110000: color_data = 12'b001110100111;
		16'b0001010010110001: color_data = 12'b001110100111;
		16'b0001010010110010: color_data = 12'b001110100111;
		16'b0001010010110011: color_data = 12'b001110100111;
		16'b0001010010110100: color_data = 12'b001110100111;
		16'b0001010010110101: color_data = 12'b001110100111;
		16'b0001010010110110: color_data = 12'b001110100111;
		16'b0001010010110111: color_data = 12'b001110100111;
		16'b0001010010111000: color_data = 12'b001110100111;
		16'b0001010010111001: color_data = 12'b001110100111;
		16'b0001010010111010: color_data = 12'b001110100111;
		16'b0001010010111011: color_data = 12'b001110100111;
		16'b0001010010111100: color_data = 12'b001110100111;
		16'b0001010010111101: color_data = 12'b001110100111;
		16'b0001010010111110: color_data = 12'b001110100111;
		16'b0001010010111111: color_data = 12'b001110100111;
		16'b0001010011000000: color_data = 12'b001110100111;
		16'b0001010011000001: color_data = 12'b001110100111;
		16'b0001010011000010: color_data = 12'b001110100111;
		16'b0001010011000011: color_data = 12'b001110100111;
		16'b0001010011000100: color_data = 12'b001110100111;
		16'b0001010011001011: color_data = 12'b001110100111;
		16'b0001010011001100: color_data = 12'b001110100111;
		16'b0001010011001101: color_data = 12'b001110100111;
		16'b0001010011001110: color_data = 12'b001110100111;
		16'b0001010011001111: color_data = 12'b001110100111;
		16'b0001010011010000: color_data = 12'b001110100111;
		16'b0001010011010001: color_data = 12'b001110100111;
		16'b0001010011010010: color_data = 12'b001110100111;
		16'b0001010011010011: color_data = 12'b001110100111;
		16'b0001010011010100: color_data = 12'b001110100111;
		16'b0001010011010101: color_data = 12'b001110100111;
		16'b0001010011010110: color_data = 12'b001110100111;
		16'b0001010011010111: color_data = 12'b001110100111;
		16'b0001010011011000: color_data = 12'b001110100111;
		16'b0001010011011001: color_data = 12'b001110100111;
		16'b0001010011011010: color_data = 12'b001110100111;
		16'b0001010011011011: color_data = 12'b001110100111;
		16'b0001010011011100: color_data = 12'b001110100111;
		16'b0001010011011101: color_data = 12'b001110100111;
		16'b0001010011011110: color_data = 12'b001110100111;
		16'b0001010011011111: color_data = 12'b001110100111;
		16'b0001010011100000: color_data = 12'b001110100111;
		16'b0001010011100001: color_data = 12'b001110100111;
		16'b0001010011100010: color_data = 12'b001110100111;
		16'b0001010011100011: color_data = 12'b001110100111;
		16'b0001010011100100: color_data = 12'b001110100111;
		16'b0001010011100101: color_data = 12'b001110100111;
		16'b0001010011100110: color_data = 12'b001110100111;
		16'b0001010011100111: color_data = 12'b001110100111;
		16'b0001010011101000: color_data = 12'b001110100111;
		16'b0001010011101001: color_data = 12'b001110100111;
		16'b0001010011101010: color_data = 12'b001110100111;
		16'b0001010011101011: color_data = 12'b001110100111;
		16'b0001010011101100: color_data = 12'b001110100111;
		16'b0001010011101101: color_data = 12'b001110100111;
		16'b0001010011101110: color_data = 12'b001110100111;
		16'b0001010011101111: color_data = 12'b001110100111;
		16'b0001010011111100: color_data = 12'b001110100111;
		16'b0001010011111101: color_data = 12'b001110100111;
		16'b0001010011111110: color_data = 12'b001110100111;
		16'b0001010011111111: color_data = 12'b001110100111;
		16'b0001010100000000: color_data = 12'b001110100111;
		16'b0001010100000001: color_data = 12'b001110100111;
		16'b0001010100000010: color_data = 12'b001110100111;
		16'b0001010100000011: color_data = 12'b001110100111;
		16'b0001010100000100: color_data = 12'b001110100111;
		16'b0001010100000101: color_data = 12'b001110100111;
		16'b0001010100000110: color_data = 12'b001110100111;
		16'b0001010100000111: color_data = 12'b001110100111;
		16'b0001010100001000: color_data = 12'b001110100111;
		16'b0001010100001001: color_data = 12'b001110100111;
		16'b0001010100001010: color_data = 12'b001110100111;
		16'b0001010100001011: color_data = 12'b001110100111;
		16'b0001010100001100: color_data = 12'b001110100111;
		16'b0001010100001101: color_data = 12'b001110100111;
		16'b0001010100001110: color_data = 12'b001110100111;
		16'b0001010100001111: color_data = 12'b001110100111;
		16'b0001010100010000: color_data = 12'b001110100111;
		16'b0001010100010001: color_data = 12'b001110100111;
		16'b0001010100010010: color_data = 12'b001110100111;
		16'b0001010100010011: color_data = 12'b001110100111;
		16'b0001010100010100: color_data = 12'b001110100111;
		16'b0001010100010101: color_data = 12'b001110100111;
		16'b0001010100010110: color_data = 12'b001110100111;
		16'b0001010100010111: color_data = 12'b001110100111;
		16'b0001010100011000: color_data = 12'b001110100111;
		16'b0001010100011001: color_data = 12'b001110100111;
		16'b0001010100011010: color_data = 12'b001110100111;
		16'b0001010100011011: color_data = 12'b001110100111;
		16'b0001010100011100: color_data = 12'b001110100111;
		16'b0001010100011101: color_data = 12'b001110100111;
		16'b0001010100011110: color_data = 12'b001110100111;
		16'b0001010100011111: color_data = 12'b001110100111;
		16'b0001010100100000: color_data = 12'b001110100111;
		16'b0001010100101101: color_data = 12'b001110100111;
		16'b0001010100101110: color_data = 12'b001110100111;
		16'b0001010100101111: color_data = 12'b001110100111;
		16'b0001010100110000: color_data = 12'b001110100111;
		16'b0001010100110001: color_data = 12'b001110100111;
		16'b0001010100110010: color_data = 12'b001110100111;
		16'b0001010100110011: color_data = 12'b001110100111;
		16'b0001010100110100: color_data = 12'b001110100111;
		16'b0001010100110101: color_data = 12'b001110100111;
		16'b0001010100110110: color_data = 12'b001110100111;
		16'b0001010100110111: color_data = 12'b001110100111;
		16'b0001010100111000: color_data = 12'b001110100111;
		16'b0001010100111001: color_data = 12'b001110100111;
		16'b0001010100111010: color_data = 12'b001110100111;
		16'b0001010100111011: color_data = 12'b001110100111;
		16'b0001010100111100: color_data = 12'b001110100111;
		16'b0001010100111101: color_data = 12'b001110100111;
		16'b0001010100111110: color_data = 12'b001110100111;
		16'b0001010100111111: color_data = 12'b001110100111;
		16'b0001010101000000: color_data = 12'b001110100111;
		16'b0001010101000001: color_data = 12'b001110100111;
		16'b0001010101000010: color_data = 12'b001110100111;
		16'b0001010101000011: color_data = 12'b001110100111;
		16'b0001010101000100: color_data = 12'b001110100111;
		16'b0001010101100100: color_data = 12'b001110100111;
		16'b0001010101100101: color_data = 12'b001110100111;
		16'b0001010101100110: color_data = 12'b001110100111;
		16'b0001010101100111: color_data = 12'b001110100111;
		16'b0001010101101000: color_data = 12'b001110100111;
		16'b0001010101101001: color_data = 12'b001110100111;
		16'b0001010101101010: color_data = 12'b001110100111;
		16'b0001010101101011: color_data = 12'b001110100111;
		16'b0001010101101100: color_data = 12'b001110100111;
		16'b0001010101101101: color_data = 12'b001110100111;
		16'b0001010101101110: color_data = 12'b001110100111;
		16'b0001010101101111: color_data = 12'b001110100111;
		16'b0001010101110000: color_data = 12'b001110100111;
		16'b0001010101110001: color_data = 12'b001110100111;
		16'b0001010101110010: color_data = 12'b001110100111;
		16'b0001010101110011: color_data = 12'b001110100111;
		16'b0001010101110100: color_data = 12'b001110100111;
		16'b0001010101110101: color_data = 12'b001110100111;
		16'b0001010101110110: color_data = 12'b001110100111;
		16'b0001010101110111: color_data = 12'b001110100111;
		16'b0001010101111000: color_data = 12'b001110100111;
		16'b0001010101111001: color_data = 12'b001110100111;
		16'b0001010101111010: color_data = 12'b001110100111;
		16'b0001010101111011: color_data = 12'b001110100111;
		16'b0001011000001101: color_data = 12'b001110100111;
		16'b0001011000001110: color_data = 12'b001110100111;
		16'b0001011000001111: color_data = 12'b001110100111;
		16'b0001011000010000: color_data = 12'b001110100111;
		16'b0001011000010001: color_data = 12'b001110100111;
		16'b0001011000010010: color_data = 12'b001110100111;
		16'b0001011000010011: color_data = 12'b001110100111;
		16'b0001011000010100: color_data = 12'b001110100111;
		16'b0001011000010101: color_data = 12'b001110100111;
		16'b0001011000010110: color_data = 12'b001110100111;
		16'b0001011000010111: color_data = 12'b001110100111;
		16'b0001011000011000: color_data = 12'b001110100111;
		16'b0001011000011001: color_data = 12'b001110100111;
		16'b0001011000011010: color_data = 12'b001110100111;
		16'b0001011000011011: color_data = 12'b001110100111;
		16'b0001011000011100: color_data = 12'b001110100111;
		16'b0001011000011101: color_data = 12'b001110100111;
		16'b0001011000011110: color_data = 12'b001110100111;
		16'b0001011000011111: color_data = 12'b001110100111;
		16'b0001011000100000: color_data = 12'b001110100111;
		16'b0001011000100001: color_data = 12'b001110100111;
		16'b0001011000100010: color_data = 12'b001110100111;
		16'b0001011000100011: color_data = 12'b001110100111;
		16'b0001011000100100: color_data = 12'b001110100111;
		16'b0001011000101011: color_data = 12'b001110100111;
		16'b0001011000101100: color_data = 12'b001110100111;
		16'b0001011000101101: color_data = 12'b001110100111;
		16'b0001011000101110: color_data = 12'b001110100111;
		16'b0001011000101111: color_data = 12'b001110100111;
		16'b0001011000110000: color_data = 12'b001110100111;
		16'b0001011000110001: color_data = 12'b001110100111;
		16'b0001011000110010: color_data = 12'b001110100111;
		16'b0001011000110011: color_data = 12'b001110100111;
		16'b0001011000110100: color_data = 12'b001110100111;
		16'b0001011000110101: color_data = 12'b001110100111;
		16'b0001011000110110: color_data = 12'b001110100111;
		16'b0001011000110111: color_data = 12'b001110100111;
		16'b0001011001000100: color_data = 12'b001110100111;
		16'b0001011001000101: color_data = 12'b001110100111;
		16'b0001011001000110: color_data = 12'b001110100111;
		16'b0001011001000111: color_data = 12'b001110100111;
		16'b0001011001001000: color_data = 12'b001110100111;
		16'b0001011001001001: color_data = 12'b001110100111;
		16'b0001011001001010: color_data = 12'b001110100111;
		16'b0001011001001011: color_data = 12'b001110100111;
		16'b0001011001001100: color_data = 12'b001110100111;
		16'b0001011001001101: color_data = 12'b001110100111;
		16'b0001011001001110: color_data = 12'b001110100111;
		16'b0001011001001111: color_data = 12'b001110100111;
		16'b0001011001010110: color_data = 12'b001110100111;
		16'b0001011001010111: color_data = 12'b001110100111;
		16'b0001011001011000: color_data = 12'b001110100111;
		16'b0001011001011001: color_data = 12'b001110100111;
		16'b0001011001011010: color_data = 12'b001110100111;
		16'b0001011001011011: color_data = 12'b001110100111;
		16'b0001011001011100: color_data = 12'b001110100111;
		16'b0001011001011101: color_data = 12'b001110100111;
		16'b0001011001011110: color_data = 12'b001110100111;
		16'b0001011001011111: color_data = 12'b001110100111;
		16'b0001011001100000: color_data = 12'b001110100111;
		16'b0001011001100001: color_data = 12'b001110100111;
		16'b0001011001100010: color_data = 12'b001110100111;
		16'b0001011001100011: color_data = 12'b001110100111;
		16'b0001011001100100: color_data = 12'b001110100111;
		16'b0001011001100101: color_data = 12'b001110100111;
		16'b0001011001100110: color_data = 12'b001110100111;
		16'b0001011001100111: color_data = 12'b001110100111;
		16'b0001011001101000: color_data = 12'b001110100111;
		16'b0001011001101001: color_data = 12'b001110100111;
		16'b0001011001101010: color_data = 12'b001110100111;
		16'b0001011001101011: color_data = 12'b001110100111;
		16'b0001011001101100: color_data = 12'b001110100111;
		16'b0001011001101101: color_data = 12'b001110100111;
		16'b0001011001101110: color_data = 12'b001110100111;
		16'b0001011001110101: color_data = 12'b001110100111;
		16'b0001011001110110: color_data = 12'b001110100111;
		16'b0001011001110111: color_data = 12'b001110100111;
		16'b0001011001111000: color_data = 12'b001110100111;
		16'b0001011001111001: color_data = 12'b001110100111;
		16'b0001011001111010: color_data = 12'b001110100111;
		16'b0001011001111011: color_data = 12'b001110100111;
		16'b0001011001111100: color_data = 12'b001110100111;
		16'b0001011001111101: color_data = 12'b001110100111;
		16'b0001011001111110: color_data = 12'b001110100111;
		16'b0001011001111111: color_data = 12'b001110100111;
		16'b0001011010000000: color_data = 12'b001110100111;
		16'b0001011010000001: color_data = 12'b001110100111;
		16'b0001011010000010: color_data = 12'b001110100111;
		16'b0001011010000011: color_data = 12'b001110100111;
		16'b0001011010000100: color_data = 12'b001110100111;
		16'b0001011010000101: color_data = 12'b001110100111;
		16'b0001011010000110: color_data = 12'b001110100111;
		16'b0001011010000111: color_data = 12'b001110100111;
		16'b0001011010001000: color_data = 12'b001110100111;
		16'b0001011010001001: color_data = 12'b001110100111;
		16'b0001011010001010: color_data = 12'b001110100111;
		16'b0001011010001011: color_data = 12'b001110100111;
		16'b0001011010001100: color_data = 12'b001110100111;
		16'b0001011010101100: color_data = 12'b001110100111;
		16'b0001011010101101: color_data = 12'b001110100111;
		16'b0001011010101110: color_data = 12'b001110100111;
		16'b0001011010101111: color_data = 12'b001110100111;
		16'b0001011010110000: color_data = 12'b001110100111;
		16'b0001011010110001: color_data = 12'b001110100111;
		16'b0001011010110010: color_data = 12'b001110100111;
		16'b0001011010110011: color_data = 12'b001110100111;
		16'b0001011010110100: color_data = 12'b001110100111;
		16'b0001011010110101: color_data = 12'b001110100111;
		16'b0001011010110110: color_data = 12'b001110100111;
		16'b0001011010110111: color_data = 12'b001110100111;
		16'b0001011010111000: color_data = 12'b001110100111;
		16'b0001011010111001: color_data = 12'b001110100111;
		16'b0001011010111010: color_data = 12'b001110100111;
		16'b0001011010111011: color_data = 12'b001110100111;
		16'b0001011010111100: color_data = 12'b001110100111;
		16'b0001011010111101: color_data = 12'b001110100111;
		16'b0001011010111110: color_data = 12'b001110100111;
		16'b0001011010111111: color_data = 12'b001110100111;
		16'b0001011011000000: color_data = 12'b001110100111;
		16'b0001011011000001: color_data = 12'b001110100111;
		16'b0001011011000010: color_data = 12'b001110100111;
		16'b0001011011000011: color_data = 12'b001110100111;
		16'b0001011011000100: color_data = 12'b001110100111;
		16'b0001011011001011: color_data = 12'b001110100111;
		16'b0001011011001100: color_data = 12'b001110100111;
		16'b0001011011001101: color_data = 12'b001110100111;
		16'b0001011011001110: color_data = 12'b001110100111;
		16'b0001011011001111: color_data = 12'b001110100111;
		16'b0001011011010000: color_data = 12'b001110100111;
		16'b0001011011010001: color_data = 12'b001110100111;
		16'b0001011011010010: color_data = 12'b001110100111;
		16'b0001011011010011: color_data = 12'b001110100111;
		16'b0001011011010100: color_data = 12'b001110100111;
		16'b0001011011010101: color_data = 12'b001110100111;
		16'b0001011011010110: color_data = 12'b001110100111;
		16'b0001011011010111: color_data = 12'b001110100111;
		16'b0001011011011000: color_data = 12'b001110100111;
		16'b0001011011011001: color_data = 12'b001110100111;
		16'b0001011011011010: color_data = 12'b001110100111;
		16'b0001011011011011: color_data = 12'b001110100111;
		16'b0001011011011100: color_data = 12'b001110100111;
		16'b0001011011011101: color_data = 12'b001110100111;
		16'b0001011011011110: color_data = 12'b001110100111;
		16'b0001011011011111: color_data = 12'b001110100111;
		16'b0001011011100000: color_data = 12'b001110100111;
		16'b0001011011100001: color_data = 12'b001110100111;
		16'b0001011011100010: color_data = 12'b001110100111;
		16'b0001011011100011: color_data = 12'b001110100111;
		16'b0001011011100100: color_data = 12'b001110100111;
		16'b0001011011100101: color_data = 12'b001110100111;
		16'b0001011011100110: color_data = 12'b001110100111;
		16'b0001011011100111: color_data = 12'b001110100111;
		16'b0001011011101000: color_data = 12'b001110100111;
		16'b0001011011101001: color_data = 12'b001110100111;
		16'b0001011011101010: color_data = 12'b001110100111;
		16'b0001011011101011: color_data = 12'b001110100111;
		16'b0001011011101100: color_data = 12'b001110100111;
		16'b0001011011101101: color_data = 12'b001110100111;
		16'b0001011011101110: color_data = 12'b001110100111;
		16'b0001011011101111: color_data = 12'b001110100111;
		16'b0001011011111100: color_data = 12'b001110100111;
		16'b0001011011111101: color_data = 12'b001110100111;
		16'b0001011011111110: color_data = 12'b001110100111;
		16'b0001011011111111: color_data = 12'b001110100111;
		16'b0001011100000000: color_data = 12'b001110100111;
		16'b0001011100000001: color_data = 12'b001110100111;
		16'b0001011100000010: color_data = 12'b001110100111;
		16'b0001011100000011: color_data = 12'b001110100111;
		16'b0001011100000100: color_data = 12'b001110100111;
		16'b0001011100000101: color_data = 12'b001110100111;
		16'b0001011100000110: color_data = 12'b001110100111;
		16'b0001011100000111: color_data = 12'b001110100111;
		16'b0001011100001000: color_data = 12'b001110100111;
		16'b0001011100001001: color_data = 12'b001110100111;
		16'b0001011100001010: color_data = 12'b001110100111;
		16'b0001011100001011: color_data = 12'b001110100111;
		16'b0001011100001100: color_data = 12'b001110100111;
		16'b0001011100001101: color_data = 12'b001110100111;
		16'b0001011100001110: color_data = 12'b001110100111;
		16'b0001011100001111: color_data = 12'b001110100111;
		16'b0001011100010000: color_data = 12'b001110100111;
		16'b0001011100010001: color_data = 12'b001110100111;
		16'b0001011100010010: color_data = 12'b001110100111;
		16'b0001011100010011: color_data = 12'b001110100111;
		16'b0001011100010100: color_data = 12'b001110100111;
		16'b0001011100010101: color_data = 12'b001110100111;
		16'b0001011100010110: color_data = 12'b001110100111;
		16'b0001011100010111: color_data = 12'b001110100111;
		16'b0001011100011000: color_data = 12'b001110100111;
		16'b0001011100011001: color_data = 12'b001110100111;
		16'b0001011100011010: color_data = 12'b001110100111;
		16'b0001011100011011: color_data = 12'b001110100111;
		16'b0001011100011100: color_data = 12'b001110100111;
		16'b0001011100011101: color_data = 12'b001110100111;
		16'b0001011100011110: color_data = 12'b001110100111;
		16'b0001011100011111: color_data = 12'b001110100111;
		16'b0001011100100000: color_data = 12'b001110100111;
		16'b0001011100101101: color_data = 12'b001110100111;
		16'b0001011100101110: color_data = 12'b001110100111;
		16'b0001011100101111: color_data = 12'b001110100111;
		16'b0001011100110000: color_data = 12'b001110100111;
		16'b0001011100110001: color_data = 12'b001110100111;
		16'b0001011100110010: color_data = 12'b001110100111;
		16'b0001011100110011: color_data = 12'b001110100111;
		16'b0001011100110100: color_data = 12'b001110100111;
		16'b0001011100110101: color_data = 12'b001110100111;
		16'b0001011100110110: color_data = 12'b001110100111;
		16'b0001011100110111: color_data = 12'b001110100111;
		16'b0001011100111000: color_data = 12'b001110100111;
		16'b0001011100111001: color_data = 12'b001110100111;
		16'b0001011100111010: color_data = 12'b001110100111;
		16'b0001011100111011: color_data = 12'b001110100111;
		16'b0001011100111100: color_data = 12'b001110100111;
		16'b0001011100111101: color_data = 12'b001110100111;
		16'b0001011100111110: color_data = 12'b001110100111;
		16'b0001011100111111: color_data = 12'b001110100111;
		16'b0001011101000000: color_data = 12'b001110100111;
		16'b0001011101000001: color_data = 12'b001110100111;
		16'b0001011101000010: color_data = 12'b001110100111;
		16'b0001011101000011: color_data = 12'b001110100111;
		16'b0001011101000100: color_data = 12'b001110100111;
		16'b0001011101100100: color_data = 12'b001110100111;
		16'b0001011101100101: color_data = 12'b001110100111;
		16'b0001011101100110: color_data = 12'b001110100111;
		16'b0001011101100111: color_data = 12'b001110100111;
		16'b0001011101101000: color_data = 12'b001110100111;
		16'b0001011101101001: color_data = 12'b001110100111;
		16'b0001011101101010: color_data = 12'b001110100111;
		16'b0001011101101011: color_data = 12'b001110100111;
		16'b0001011101101100: color_data = 12'b001110100111;
		16'b0001011101101101: color_data = 12'b001110100111;
		16'b0001011101101110: color_data = 12'b001110100111;
		16'b0001011101101111: color_data = 12'b001110100111;
		16'b0001011101110000: color_data = 12'b001110100111;
		16'b0001011101110001: color_data = 12'b001110100111;
		16'b0001011101110010: color_data = 12'b001110100111;
		16'b0001011101110011: color_data = 12'b001110100111;
		16'b0001011101110100: color_data = 12'b001110100111;
		16'b0001011101110101: color_data = 12'b001110100111;
		16'b0001011101110110: color_data = 12'b001110100111;
		16'b0001011101110111: color_data = 12'b001110100111;
		16'b0001011101111000: color_data = 12'b001110100111;
		16'b0001011101111001: color_data = 12'b001110100111;
		16'b0001011101111010: color_data = 12'b001110100111;
		16'b0001011101111011: color_data = 12'b001110100111;
		16'b0001100000001101: color_data = 12'b001110100111;
		16'b0001100000001110: color_data = 12'b001110100111;
		16'b0001100000001111: color_data = 12'b001110100111;
		16'b0001100000010000: color_data = 12'b001110100111;
		16'b0001100000010001: color_data = 12'b001110100111;
		16'b0001100000010010: color_data = 12'b001110100111;
		16'b0001100000010011: color_data = 12'b001110100111;
		16'b0001100000010100: color_data = 12'b001110100111;
		16'b0001100000010101: color_data = 12'b001110100111;
		16'b0001100000010110: color_data = 12'b001110100111;
		16'b0001100000010111: color_data = 12'b001110100111;
		16'b0001100000011000: color_data = 12'b001110100111;
		16'b0001100000011001: color_data = 12'b001110100111;
		16'b0001100000011010: color_data = 12'b001110100111;
		16'b0001100000011011: color_data = 12'b001110100111;
		16'b0001100000011100: color_data = 12'b001110100111;
		16'b0001100000011101: color_data = 12'b001110100111;
		16'b0001100000011110: color_data = 12'b001110100111;
		16'b0001100000011111: color_data = 12'b001110100111;
		16'b0001100000100000: color_data = 12'b001110100111;
		16'b0001100000100001: color_data = 12'b001110100111;
		16'b0001100000100010: color_data = 12'b001110100111;
		16'b0001100000100011: color_data = 12'b001110100111;
		16'b0001100000100100: color_data = 12'b001110100111;
		16'b0001100000101011: color_data = 12'b001110100111;
		16'b0001100000101100: color_data = 12'b001110100111;
		16'b0001100000101101: color_data = 12'b001110100111;
		16'b0001100000101110: color_data = 12'b001110100111;
		16'b0001100000101111: color_data = 12'b001110100111;
		16'b0001100000110000: color_data = 12'b001110100111;
		16'b0001100000110001: color_data = 12'b001110100111;
		16'b0001100000110010: color_data = 12'b001110100111;
		16'b0001100000110011: color_data = 12'b001110100111;
		16'b0001100000110100: color_data = 12'b001110100111;
		16'b0001100000110101: color_data = 12'b001110100111;
		16'b0001100000110110: color_data = 12'b001110100111;
		16'b0001100000110111: color_data = 12'b001110100111;
		16'b0001100001000100: color_data = 12'b001110100111;
		16'b0001100001000101: color_data = 12'b001110100111;
		16'b0001100001000110: color_data = 12'b001110100111;
		16'b0001100001000111: color_data = 12'b001110100111;
		16'b0001100001001000: color_data = 12'b001110100111;
		16'b0001100001001001: color_data = 12'b001110100111;
		16'b0001100001001010: color_data = 12'b001110100111;
		16'b0001100001001011: color_data = 12'b001110100111;
		16'b0001100001001100: color_data = 12'b001110100111;
		16'b0001100001001101: color_data = 12'b001110100111;
		16'b0001100001001110: color_data = 12'b001110100111;
		16'b0001100001001111: color_data = 12'b001110100111;
		16'b0001100001010110: color_data = 12'b001110100111;
		16'b0001100001010111: color_data = 12'b001110100111;
		16'b0001100001011000: color_data = 12'b001110100111;
		16'b0001100001011001: color_data = 12'b001110100111;
		16'b0001100001011010: color_data = 12'b001110100111;
		16'b0001100001011011: color_data = 12'b001110100111;
		16'b0001100001011100: color_data = 12'b001110100111;
		16'b0001100001011101: color_data = 12'b001110100111;
		16'b0001100001011110: color_data = 12'b001110100111;
		16'b0001100001011111: color_data = 12'b001110100111;
		16'b0001100001100000: color_data = 12'b001110100111;
		16'b0001100001100001: color_data = 12'b001110100111;
		16'b0001100001100010: color_data = 12'b001110100111;
		16'b0001100001100011: color_data = 12'b001110100111;
		16'b0001100001100100: color_data = 12'b001110100111;
		16'b0001100001100101: color_data = 12'b001110100111;
		16'b0001100001100110: color_data = 12'b001110100111;
		16'b0001100001100111: color_data = 12'b001110100111;
		16'b0001100001101000: color_data = 12'b001110100111;
		16'b0001100001101001: color_data = 12'b001110100111;
		16'b0001100001101010: color_data = 12'b001110100111;
		16'b0001100001101011: color_data = 12'b001110100111;
		16'b0001100001101100: color_data = 12'b001110100111;
		16'b0001100001101101: color_data = 12'b001110100111;
		16'b0001100001101110: color_data = 12'b001110100111;
		16'b0001100001110101: color_data = 12'b001110100111;
		16'b0001100001110110: color_data = 12'b001110100111;
		16'b0001100001110111: color_data = 12'b001110100111;
		16'b0001100001111000: color_data = 12'b001110100111;
		16'b0001100001111001: color_data = 12'b001110100111;
		16'b0001100001111010: color_data = 12'b001110100111;
		16'b0001100001111011: color_data = 12'b001110100111;
		16'b0001100001111100: color_data = 12'b001110100111;
		16'b0001100001111101: color_data = 12'b001110100111;
		16'b0001100001111110: color_data = 12'b001110100111;
		16'b0001100001111111: color_data = 12'b001110100111;
		16'b0001100010000000: color_data = 12'b001110100111;
		16'b0001100010000001: color_data = 12'b001110100111;
		16'b0001100010000010: color_data = 12'b001110100111;
		16'b0001100010000011: color_data = 12'b001110100111;
		16'b0001100010000100: color_data = 12'b001110100111;
		16'b0001100010000101: color_data = 12'b001110100111;
		16'b0001100010000110: color_data = 12'b001110100111;
		16'b0001100010000111: color_data = 12'b001110100111;
		16'b0001100010001000: color_data = 12'b001110100111;
		16'b0001100010001001: color_data = 12'b001110100111;
		16'b0001100010001010: color_data = 12'b001110100111;
		16'b0001100010001011: color_data = 12'b001110100111;
		16'b0001100010001100: color_data = 12'b001110100111;
		16'b0001100010101100: color_data = 12'b001110100111;
		16'b0001100010101101: color_data = 12'b001110100111;
		16'b0001100010101110: color_data = 12'b001110100111;
		16'b0001100010101111: color_data = 12'b001110100111;
		16'b0001100010110000: color_data = 12'b001110100111;
		16'b0001100010110001: color_data = 12'b001110100111;
		16'b0001100010110010: color_data = 12'b001110100111;
		16'b0001100010110011: color_data = 12'b001110100111;
		16'b0001100010110100: color_data = 12'b001110100111;
		16'b0001100010110101: color_data = 12'b001110100111;
		16'b0001100010110110: color_data = 12'b001110100111;
		16'b0001100010110111: color_data = 12'b001110100111;
		16'b0001100010111000: color_data = 12'b001110100111;
		16'b0001100010111001: color_data = 12'b001110100111;
		16'b0001100010111010: color_data = 12'b001110100111;
		16'b0001100010111011: color_data = 12'b001110100111;
		16'b0001100010111100: color_data = 12'b001110100111;
		16'b0001100010111101: color_data = 12'b001110100111;
		16'b0001100010111110: color_data = 12'b001110100111;
		16'b0001100010111111: color_data = 12'b001110100111;
		16'b0001100011000000: color_data = 12'b001110100111;
		16'b0001100011000001: color_data = 12'b001110100111;
		16'b0001100011000010: color_data = 12'b001110100111;
		16'b0001100011000011: color_data = 12'b001110100111;
		16'b0001100011000100: color_data = 12'b001110100111;
		16'b0001100011001011: color_data = 12'b001110100111;
		16'b0001100011001100: color_data = 12'b001110100111;
		16'b0001100011001101: color_data = 12'b001110100111;
		16'b0001100011001110: color_data = 12'b001110100111;
		16'b0001100011001111: color_data = 12'b001110100111;
		16'b0001100011010000: color_data = 12'b001110100111;
		16'b0001100011010001: color_data = 12'b001110100111;
		16'b0001100011010010: color_data = 12'b001110100111;
		16'b0001100011010011: color_data = 12'b001110100111;
		16'b0001100011010100: color_data = 12'b001110100111;
		16'b0001100011010101: color_data = 12'b001110100111;
		16'b0001100011010110: color_data = 12'b001110100111;
		16'b0001100011010111: color_data = 12'b001110100111;
		16'b0001100011011000: color_data = 12'b001110100111;
		16'b0001100011011001: color_data = 12'b001110100111;
		16'b0001100011011010: color_data = 12'b001110100111;
		16'b0001100011011011: color_data = 12'b001110100111;
		16'b0001100011011100: color_data = 12'b001110100111;
		16'b0001100011011101: color_data = 12'b001110100111;
		16'b0001100011011110: color_data = 12'b001110100111;
		16'b0001100011011111: color_data = 12'b001110100111;
		16'b0001100011100000: color_data = 12'b001110100111;
		16'b0001100011100001: color_data = 12'b001110100111;
		16'b0001100011100010: color_data = 12'b001110100111;
		16'b0001100011100011: color_data = 12'b001110100111;
		16'b0001100011100100: color_data = 12'b001110100111;
		16'b0001100011100101: color_data = 12'b001110100111;
		16'b0001100011100110: color_data = 12'b001110100111;
		16'b0001100011100111: color_data = 12'b001110100111;
		16'b0001100011101000: color_data = 12'b001110100111;
		16'b0001100011101001: color_data = 12'b001110100111;
		16'b0001100011101010: color_data = 12'b001110100111;
		16'b0001100011101011: color_data = 12'b001110100111;
		16'b0001100011101100: color_data = 12'b001110100111;
		16'b0001100011101101: color_data = 12'b001110100111;
		16'b0001100011101110: color_data = 12'b001110100111;
		16'b0001100011101111: color_data = 12'b001110100111;
		16'b0001100011111100: color_data = 12'b001110100111;
		16'b0001100011111101: color_data = 12'b001110100111;
		16'b0001100011111110: color_data = 12'b001110100111;
		16'b0001100011111111: color_data = 12'b001110100111;
		16'b0001100100000000: color_data = 12'b001110100111;
		16'b0001100100000001: color_data = 12'b001110100111;
		16'b0001100100000010: color_data = 12'b001110100111;
		16'b0001100100000011: color_data = 12'b001110100111;
		16'b0001100100000100: color_data = 12'b001110100111;
		16'b0001100100000101: color_data = 12'b001110100111;
		16'b0001100100000110: color_data = 12'b001110100111;
		16'b0001100100000111: color_data = 12'b001110100111;
		16'b0001100100001000: color_data = 12'b001110100111;
		16'b0001100100001001: color_data = 12'b001110100111;
		16'b0001100100001010: color_data = 12'b001110100111;
		16'b0001100100001011: color_data = 12'b001110100111;
		16'b0001100100001100: color_data = 12'b001110100111;
		16'b0001100100001101: color_data = 12'b001110100111;
		16'b0001100100001110: color_data = 12'b001110100111;
		16'b0001100100001111: color_data = 12'b001110100111;
		16'b0001100100010000: color_data = 12'b001110100111;
		16'b0001100100010001: color_data = 12'b001110100111;
		16'b0001100100010010: color_data = 12'b001110100111;
		16'b0001100100010011: color_data = 12'b001110100111;
		16'b0001100100010100: color_data = 12'b001110100111;
		16'b0001100100010101: color_data = 12'b001110100111;
		16'b0001100100010110: color_data = 12'b001110100111;
		16'b0001100100010111: color_data = 12'b001110100111;
		16'b0001100100011000: color_data = 12'b001110100111;
		16'b0001100100011001: color_data = 12'b001110100111;
		16'b0001100100011010: color_data = 12'b001110100111;
		16'b0001100100011011: color_data = 12'b001110100111;
		16'b0001100100011100: color_data = 12'b001110100111;
		16'b0001100100011101: color_data = 12'b001110100111;
		16'b0001100100011110: color_data = 12'b001110100111;
		16'b0001100100011111: color_data = 12'b001110100111;
		16'b0001100100100000: color_data = 12'b001110100111;
		16'b0001100100101101: color_data = 12'b001110100111;
		16'b0001100100101110: color_data = 12'b001110100111;
		16'b0001100100101111: color_data = 12'b001110100111;
		16'b0001100100110000: color_data = 12'b001110100111;
		16'b0001100100110001: color_data = 12'b001110100111;
		16'b0001100100110010: color_data = 12'b001110100111;
		16'b0001100100110011: color_data = 12'b001110100111;
		16'b0001100100110100: color_data = 12'b001110100111;
		16'b0001100100110101: color_data = 12'b001110100111;
		16'b0001100100110110: color_data = 12'b001110100111;
		16'b0001100100110111: color_data = 12'b001110100111;
		16'b0001100100111000: color_data = 12'b001110100111;
		16'b0001100100111001: color_data = 12'b001110100111;
		16'b0001100100111010: color_data = 12'b001110100111;
		16'b0001100100111011: color_data = 12'b001110100111;
		16'b0001100100111100: color_data = 12'b001110100111;
		16'b0001100100111101: color_data = 12'b001110100111;
		16'b0001100100111110: color_data = 12'b001110100111;
		16'b0001100100111111: color_data = 12'b001110100111;
		16'b0001100101000000: color_data = 12'b001110100111;
		16'b0001100101000001: color_data = 12'b001110100111;
		16'b0001100101000010: color_data = 12'b001110100111;
		16'b0001100101000011: color_data = 12'b001110100111;
		16'b0001100101000100: color_data = 12'b001110100111;
		16'b0001100101100100: color_data = 12'b001110100111;
		16'b0001100101100101: color_data = 12'b001110100111;
		16'b0001100101100110: color_data = 12'b001110100111;
		16'b0001100101100111: color_data = 12'b001110100111;
		16'b0001100101101000: color_data = 12'b001110100111;
		16'b0001100101101001: color_data = 12'b001110100111;
		16'b0001100101101010: color_data = 12'b001110100111;
		16'b0001100101101011: color_data = 12'b001110100111;
		16'b0001100101101100: color_data = 12'b001110100111;
		16'b0001100101101101: color_data = 12'b001110100111;
		16'b0001100101101110: color_data = 12'b001110100111;
		16'b0001100101101111: color_data = 12'b001110100111;
		16'b0001100101110000: color_data = 12'b001110100111;
		16'b0001100101110001: color_data = 12'b001110100111;
		16'b0001100101110010: color_data = 12'b001110100111;
		16'b0001100101110011: color_data = 12'b001110100111;
		16'b0001100101110100: color_data = 12'b001110100111;
		16'b0001100101110101: color_data = 12'b001110100111;
		16'b0001100101110110: color_data = 12'b001110100111;
		16'b0001100101110111: color_data = 12'b001110100111;
		16'b0001100101111000: color_data = 12'b001110100111;
		16'b0001100101111001: color_data = 12'b001110100111;
		16'b0001100101111010: color_data = 12'b001110100111;
		16'b0001100101111011: color_data = 12'b001110100111;
		16'b0001101000000111: color_data = 12'b001110100111;
		16'b0001101000001000: color_data = 12'b001110100111;
		16'b0001101000001001: color_data = 12'b001110100111;
		16'b0001101000001010: color_data = 12'b001110100111;
		16'b0001101000001011: color_data = 12'b001110100111;
		16'b0001101000001100: color_data = 12'b001110100111;
		16'b0001101000001101: color_data = 12'b001110100111;
		16'b0001101000001110: color_data = 12'b001110100111;
		16'b0001101000001111: color_data = 12'b001110100111;
		16'b0001101000010000: color_data = 12'b001110100111;
		16'b0001101000010001: color_data = 12'b001110100111;
		16'b0001101000010010: color_data = 12'b001110100111;
		16'b0001101000010011: color_data = 12'b001110100111;
		16'b0001101000010100: color_data = 12'b001110100111;
		16'b0001101000010101: color_data = 12'b001110100111;
		16'b0001101000010110: color_data = 12'b001110100111;
		16'b0001101000010111: color_data = 12'b001110100111;
		16'b0001101000011000: color_data = 12'b001110100111;
		16'b0001101000011001: color_data = 12'b001110100111;
		16'b0001101000011010: color_data = 12'b001110100111;
		16'b0001101000011011: color_data = 12'b001110100111;
		16'b0001101000011100: color_data = 12'b001110100111;
		16'b0001101000011101: color_data = 12'b001110100111;
		16'b0001101000011110: color_data = 12'b001110100111;
		16'b0001101000011111: color_data = 12'b001110100111;
		16'b0001101000100000: color_data = 12'b001110100111;
		16'b0001101000100001: color_data = 12'b001110100111;
		16'b0001101000100010: color_data = 12'b001110100111;
		16'b0001101000100011: color_data = 12'b001110100111;
		16'b0001101000100100: color_data = 12'b001110100111;
		16'b0001101000101011: color_data = 12'b001110100111;
		16'b0001101000101100: color_data = 12'b001110100111;
		16'b0001101000101101: color_data = 12'b001110100111;
		16'b0001101000101110: color_data = 12'b001110100111;
		16'b0001101000101111: color_data = 12'b001110100111;
		16'b0001101000110000: color_data = 12'b001110100111;
		16'b0001101000110001: color_data = 12'b001110100111;
		16'b0001101000110010: color_data = 12'b001110100111;
		16'b0001101000110011: color_data = 12'b001110100111;
		16'b0001101000110100: color_data = 12'b001110100111;
		16'b0001101000110101: color_data = 12'b001110100111;
		16'b0001101000110110: color_data = 12'b001110100111;
		16'b0001101000110111: color_data = 12'b001110100111;
		16'b0001101001000100: color_data = 12'b001110100111;
		16'b0001101001000101: color_data = 12'b001110100111;
		16'b0001101001000110: color_data = 12'b001110100111;
		16'b0001101001000111: color_data = 12'b001110100111;
		16'b0001101001001000: color_data = 12'b001110100111;
		16'b0001101001001001: color_data = 12'b001110100111;
		16'b0001101001001010: color_data = 12'b001110100111;
		16'b0001101001001011: color_data = 12'b001110100111;
		16'b0001101001001100: color_data = 12'b001110100111;
		16'b0001101001001101: color_data = 12'b001110100111;
		16'b0001101001001110: color_data = 12'b001110100111;
		16'b0001101001001111: color_data = 12'b001110100111;
		16'b0001101001010110: color_data = 12'b001110100111;
		16'b0001101001010111: color_data = 12'b001110100111;
		16'b0001101001011000: color_data = 12'b001110100111;
		16'b0001101001011001: color_data = 12'b001110100111;
		16'b0001101001011010: color_data = 12'b001110100111;
		16'b0001101001011011: color_data = 12'b001110100111;
		16'b0001101001011100: color_data = 12'b001110100111;
		16'b0001101001011101: color_data = 12'b001110100111;
		16'b0001101001011110: color_data = 12'b001110100111;
		16'b0001101001011111: color_data = 12'b001110100111;
		16'b0001101001100000: color_data = 12'b001110100111;
		16'b0001101001100001: color_data = 12'b001110100111;
		16'b0001101001100010: color_data = 12'b001110100111;
		16'b0001101001100011: color_data = 12'b001110100111;
		16'b0001101001100100: color_data = 12'b001110100111;
		16'b0001101001100101: color_data = 12'b001110100111;
		16'b0001101001100110: color_data = 12'b001110100111;
		16'b0001101001100111: color_data = 12'b001110100111;
		16'b0001101001101000: color_data = 12'b001110100111;
		16'b0001101001101001: color_data = 12'b001110100111;
		16'b0001101001101010: color_data = 12'b001110100111;
		16'b0001101001101011: color_data = 12'b001110100111;
		16'b0001101001101100: color_data = 12'b001110100111;
		16'b0001101001101101: color_data = 12'b001110100111;
		16'b0001101001101110: color_data = 12'b001110100111;
		16'b0001101001110101: color_data = 12'b001110100111;
		16'b0001101001110110: color_data = 12'b001110100111;
		16'b0001101001110111: color_data = 12'b001110100111;
		16'b0001101001111000: color_data = 12'b001110100111;
		16'b0001101001111001: color_data = 12'b001110100111;
		16'b0001101001111010: color_data = 12'b001110100111;
		16'b0001101001111011: color_data = 12'b001110100111;
		16'b0001101001111100: color_data = 12'b001110100111;
		16'b0001101001111101: color_data = 12'b001110100111;
		16'b0001101001111110: color_data = 12'b001110100111;
		16'b0001101001111111: color_data = 12'b001110100111;
		16'b0001101010000000: color_data = 12'b001110100111;
		16'b0001101010000001: color_data = 12'b001110100111;
		16'b0001101010000010: color_data = 12'b001110100111;
		16'b0001101010000011: color_data = 12'b001110100111;
		16'b0001101010000100: color_data = 12'b001110100111;
		16'b0001101010000101: color_data = 12'b001110100111;
		16'b0001101010000110: color_data = 12'b001110100111;
		16'b0001101010000111: color_data = 12'b001110100111;
		16'b0001101010001000: color_data = 12'b001110100111;
		16'b0001101010001001: color_data = 12'b001110100111;
		16'b0001101010001010: color_data = 12'b001110100111;
		16'b0001101010001011: color_data = 12'b001110100111;
		16'b0001101010001100: color_data = 12'b001110100111;
		16'b0001101010001101: color_data = 12'b001110100111;
		16'b0001101010001110: color_data = 12'b001110100111;
		16'b0001101010001111: color_data = 12'b001110100111;
		16'b0001101010010000: color_data = 12'b001110100111;
		16'b0001101010010001: color_data = 12'b001110100111;
		16'b0001101010010010: color_data = 12'b001110100111;
		16'b0001101010010011: color_data = 12'b001110100111;
		16'b0001101010100110: color_data = 12'b001110100111;
		16'b0001101010100111: color_data = 12'b001110100111;
		16'b0001101010101000: color_data = 12'b001110100111;
		16'b0001101010101001: color_data = 12'b001110100111;
		16'b0001101010101010: color_data = 12'b001110100111;
		16'b0001101010101011: color_data = 12'b001110100111;
		16'b0001101010101100: color_data = 12'b001110100111;
		16'b0001101010101101: color_data = 12'b001110100111;
		16'b0001101010101110: color_data = 12'b001110100111;
		16'b0001101010101111: color_data = 12'b001110100111;
		16'b0001101010110000: color_data = 12'b001110100111;
		16'b0001101010110001: color_data = 12'b001110100111;
		16'b0001101010110010: color_data = 12'b001110100111;
		16'b0001101010110011: color_data = 12'b001110100111;
		16'b0001101010110100: color_data = 12'b001110100111;
		16'b0001101010110101: color_data = 12'b001110100111;
		16'b0001101010110110: color_data = 12'b001110100111;
		16'b0001101010110111: color_data = 12'b001110100111;
		16'b0001101010111000: color_data = 12'b001110100111;
		16'b0001101010111001: color_data = 12'b001110100111;
		16'b0001101010111010: color_data = 12'b001110100111;
		16'b0001101010111011: color_data = 12'b001110100111;
		16'b0001101010111100: color_data = 12'b001110100111;
		16'b0001101010111101: color_data = 12'b001110100111;
		16'b0001101010111110: color_data = 12'b001110100111;
		16'b0001101010111111: color_data = 12'b001110100111;
		16'b0001101011000000: color_data = 12'b001110100111;
		16'b0001101011000001: color_data = 12'b001110100111;
		16'b0001101011000010: color_data = 12'b001110100111;
		16'b0001101011000011: color_data = 12'b001110100111;
		16'b0001101011000100: color_data = 12'b001110100111;
		16'b0001101011001011: color_data = 12'b001110100111;
		16'b0001101011001100: color_data = 12'b001110100111;
		16'b0001101011001101: color_data = 12'b001110100111;
		16'b0001101011001110: color_data = 12'b001110100111;
		16'b0001101011001111: color_data = 12'b001110100111;
		16'b0001101011010000: color_data = 12'b001110100111;
		16'b0001101011010001: color_data = 12'b001110100111;
		16'b0001101011010010: color_data = 12'b001110100111;
		16'b0001101011010011: color_data = 12'b001110100111;
		16'b0001101011010100: color_data = 12'b001110100111;
		16'b0001101011010101: color_data = 12'b001110100111;
		16'b0001101011010110: color_data = 12'b001110100111;
		16'b0001101011010111: color_data = 12'b001110100111;
		16'b0001101011011000: color_data = 12'b001110100111;
		16'b0001101011011001: color_data = 12'b001110100111;
		16'b0001101011011010: color_data = 12'b001110100111;
		16'b0001101011011011: color_data = 12'b001110100111;
		16'b0001101011011100: color_data = 12'b001110100111;
		16'b0001101011011101: color_data = 12'b001110100111;
		16'b0001101011011110: color_data = 12'b001110100111;
		16'b0001101011011111: color_data = 12'b001110100111;
		16'b0001101011100000: color_data = 12'b001110100111;
		16'b0001101011100001: color_data = 12'b001110100111;
		16'b0001101011100010: color_data = 12'b001110100111;
		16'b0001101011100011: color_data = 12'b001110100111;
		16'b0001101011100100: color_data = 12'b001110100111;
		16'b0001101011100101: color_data = 12'b001110100111;
		16'b0001101011100110: color_data = 12'b001110100111;
		16'b0001101011100111: color_data = 12'b001110100111;
		16'b0001101011101000: color_data = 12'b001110100111;
		16'b0001101011101001: color_data = 12'b001110100111;
		16'b0001101011101010: color_data = 12'b001110100111;
		16'b0001101011101011: color_data = 12'b001110100111;
		16'b0001101011101100: color_data = 12'b001110100111;
		16'b0001101011101101: color_data = 12'b001110100111;
		16'b0001101011101110: color_data = 12'b001110100111;
		16'b0001101011101111: color_data = 12'b001110100111;
		16'b0001101011110110: color_data = 12'b001110100111;
		16'b0001101011110111: color_data = 12'b001110100111;
		16'b0001101011111000: color_data = 12'b001110100111;
		16'b0001101011111001: color_data = 12'b001110100111;
		16'b0001101011111010: color_data = 12'b001110100111;
		16'b0001101011111011: color_data = 12'b001110100111;
		16'b0001101011111100: color_data = 12'b001110100111;
		16'b0001101011111101: color_data = 12'b001110100111;
		16'b0001101011111110: color_data = 12'b001110100111;
		16'b0001101011111111: color_data = 12'b001110100111;
		16'b0001101100000000: color_data = 12'b001110100111;
		16'b0001101100000001: color_data = 12'b001110100111;
		16'b0001101100000010: color_data = 12'b001110100111;
		16'b0001101100000011: color_data = 12'b001110100111;
		16'b0001101100000100: color_data = 12'b001110100111;
		16'b0001101100000101: color_data = 12'b001110100111;
		16'b0001101100000110: color_data = 12'b001110100111;
		16'b0001101100000111: color_data = 12'b001110100111;
		16'b0001101100001000: color_data = 12'b001110100111;
		16'b0001101100001001: color_data = 12'b001110100111;
		16'b0001101100001010: color_data = 12'b001110100111;
		16'b0001101100001011: color_data = 12'b001110100111;
		16'b0001101100001100: color_data = 12'b001110100111;
		16'b0001101100001101: color_data = 12'b001110100111;
		16'b0001101100001110: color_data = 12'b001110100111;
		16'b0001101100001111: color_data = 12'b001110100111;
		16'b0001101100010000: color_data = 12'b001110100111;
		16'b0001101100010001: color_data = 12'b001110100111;
		16'b0001101100010010: color_data = 12'b001110100111;
		16'b0001101100010011: color_data = 12'b001110100111;
		16'b0001101100010100: color_data = 12'b001110100111;
		16'b0001101100010101: color_data = 12'b001110100111;
		16'b0001101100010110: color_data = 12'b001110100111;
		16'b0001101100010111: color_data = 12'b001110100111;
		16'b0001101100011000: color_data = 12'b001110100111;
		16'b0001101100011001: color_data = 12'b001110100111;
		16'b0001101100011010: color_data = 12'b001110100111;
		16'b0001101100011011: color_data = 12'b001110100111;
		16'b0001101100011100: color_data = 12'b001110100111;
		16'b0001101100011101: color_data = 12'b001110100111;
		16'b0001101100011110: color_data = 12'b001110100111;
		16'b0001101100011111: color_data = 12'b001110100111;
		16'b0001101100100000: color_data = 12'b001110100111;
		16'b0001101100100001: color_data = 12'b001110100111;
		16'b0001101100100010: color_data = 12'b001110100111;
		16'b0001101100100011: color_data = 12'b001110100111;
		16'b0001101100100100: color_data = 12'b001110100111;
		16'b0001101100100101: color_data = 12'b001110100111;
		16'b0001101100100110: color_data = 12'b001110100111;
		16'b0001101100101101: color_data = 12'b001110100111;
		16'b0001101100101110: color_data = 12'b001110100111;
		16'b0001101100101111: color_data = 12'b001110100111;
		16'b0001101100110000: color_data = 12'b001110100111;
		16'b0001101100110001: color_data = 12'b001110100111;
		16'b0001101100110010: color_data = 12'b001110100111;
		16'b0001101100110011: color_data = 12'b001110100111;
		16'b0001101100110100: color_data = 12'b001110100111;
		16'b0001101100110101: color_data = 12'b001110100111;
		16'b0001101100110110: color_data = 12'b001110100111;
		16'b0001101100110111: color_data = 12'b001110100111;
		16'b0001101100111000: color_data = 12'b001110100111;
		16'b0001101100111001: color_data = 12'b001110100111;
		16'b0001101100111010: color_data = 12'b001110100111;
		16'b0001101100111011: color_data = 12'b001110100111;
		16'b0001101100111100: color_data = 12'b001110100111;
		16'b0001101100111101: color_data = 12'b001110100111;
		16'b0001101100111110: color_data = 12'b001110100111;
		16'b0001101100111111: color_data = 12'b001110100111;
		16'b0001101101000000: color_data = 12'b001110100111;
		16'b0001101101000001: color_data = 12'b001110100111;
		16'b0001101101000010: color_data = 12'b001110100111;
		16'b0001101101000011: color_data = 12'b001110100111;
		16'b0001101101000100: color_data = 12'b001110100111;
		16'b0001101101000101: color_data = 12'b001110100111;
		16'b0001101101000110: color_data = 12'b001110100111;
		16'b0001101101000111: color_data = 12'b001110100111;
		16'b0001101101001000: color_data = 12'b001110100111;
		16'b0001101101001001: color_data = 12'b001110100111;
		16'b0001101101001010: color_data = 12'b001110100111;
		16'b0001101101011110: color_data = 12'b001110100111;
		16'b0001101101011111: color_data = 12'b001110100111;
		16'b0001101101100000: color_data = 12'b001110100111;
		16'b0001101101100001: color_data = 12'b001110100111;
		16'b0001101101100010: color_data = 12'b001110100111;
		16'b0001101101100011: color_data = 12'b001110100111;
		16'b0001101101100100: color_data = 12'b001110100111;
		16'b0001101101100101: color_data = 12'b001110100111;
		16'b0001101101100110: color_data = 12'b001110100111;
		16'b0001101101100111: color_data = 12'b001110100111;
		16'b0001101101101000: color_data = 12'b001110100111;
		16'b0001101101101001: color_data = 12'b001110100111;
		16'b0001101101101010: color_data = 12'b001110100111;
		16'b0001101101101011: color_data = 12'b001110100111;
		16'b0001101101101100: color_data = 12'b001110100111;
		16'b0001101101101101: color_data = 12'b001110100111;
		16'b0001101101101110: color_data = 12'b001110100111;
		16'b0001101101101111: color_data = 12'b001110100111;
		16'b0001101101110000: color_data = 12'b001110100111;
		16'b0001101101110001: color_data = 12'b001110100111;
		16'b0001101101110010: color_data = 12'b001110100111;
		16'b0001101101110011: color_data = 12'b001110100111;
		16'b0001101101110100: color_data = 12'b001110100111;
		16'b0001101101110101: color_data = 12'b001110100111;
		16'b0001101101110110: color_data = 12'b001110100111;
		16'b0001101101110111: color_data = 12'b001110100111;
		16'b0001101101111000: color_data = 12'b001110100111;
		16'b0001101101111001: color_data = 12'b001110100111;
		16'b0001101101111010: color_data = 12'b001110100111;
		16'b0001101101111011: color_data = 12'b001110100111;
		16'b0001110000000111: color_data = 12'b001110100111;
		16'b0001110000001000: color_data = 12'b001110100111;
		16'b0001110000001001: color_data = 12'b001110100111;
		16'b0001110000001010: color_data = 12'b001110100111;
		16'b0001110000001011: color_data = 12'b001110100111;
		16'b0001110000001100: color_data = 12'b001110100111;
		16'b0001110000001101: color_data = 12'b001110100111;
		16'b0001110000001110: color_data = 12'b001110100111;
		16'b0001110000001111: color_data = 12'b001110100111;
		16'b0001110000010000: color_data = 12'b001110100111;
		16'b0001110000010001: color_data = 12'b001110100111;
		16'b0001110000010010: color_data = 12'b001110100111;
		16'b0001110000010011: color_data = 12'b001110100111;
		16'b0001110000010100: color_data = 12'b001110100111;
		16'b0001110000010101: color_data = 12'b001110100111;
		16'b0001110000010110: color_data = 12'b001110100111;
		16'b0001110000010111: color_data = 12'b001110100111;
		16'b0001110000011000: color_data = 12'b001110100111;
		16'b0001110000011001: color_data = 12'b001110100111;
		16'b0001110000011010: color_data = 12'b001110100111;
		16'b0001110000011011: color_data = 12'b001110100111;
		16'b0001110000011100: color_data = 12'b001110100111;
		16'b0001110000011101: color_data = 12'b001110100111;
		16'b0001110000011110: color_data = 12'b001110100111;
		16'b0001110000011111: color_data = 12'b001110100111;
		16'b0001110000100000: color_data = 12'b001110100111;
		16'b0001110000100001: color_data = 12'b001110100111;
		16'b0001110000100010: color_data = 12'b001110100111;
		16'b0001110000100011: color_data = 12'b001110100111;
		16'b0001110000100100: color_data = 12'b001110100111;
		16'b0001110000101011: color_data = 12'b001110100111;
		16'b0001110000101100: color_data = 12'b001110100111;
		16'b0001110000101101: color_data = 12'b001110100111;
		16'b0001110000101110: color_data = 12'b001110100111;
		16'b0001110000101111: color_data = 12'b001110100111;
		16'b0001110000110000: color_data = 12'b001110100111;
		16'b0001110000110001: color_data = 12'b001110100111;
		16'b0001110000110010: color_data = 12'b001110100111;
		16'b0001110000110011: color_data = 12'b001110100111;
		16'b0001110000110100: color_data = 12'b001110100111;
		16'b0001110000110101: color_data = 12'b001110100111;
		16'b0001110000110110: color_data = 12'b001110100111;
		16'b0001110000110111: color_data = 12'b001110100111;
		16'b0001110001000100: color_data = 12'b001110100111;
		16'b0001110001000101: color_data = 12'b001110100111;
		16'b0001110001000110: color_data = 12'b001110100111;
		16'b0001110001000111: color_data = 12'b001110100111;
		16'b0001110001001000: color_data = 12'b001110100111;
		16'b0001110001001001: color_data = 12'b001110100111;
		16'b0001110001001010: color_data = 12'b001110100111;
		16'b0001110001001011: color_data = 12'b001110100111;
		16'b0001110001001100: color_data = 12'b001110100111;
		16'b0001110001001101: color_data = 12'b001110100111;
		16'b0001110001001110: color_data = 12'b001110100111;
		16'b0001110001001111: color_data = 12'b001110100111;
		16'b0001110001010110: color_data = 12'b001110100111;
		16'b0001110001010111: color_data = 12'b001110100111;
		16'b0001110001011000: color_data = 12'b001110100111;
		16'b0001110001011001: color_data = 12'b001110100111;
		16'b0001110001011010: color_data = 12'b001110100111;
		16'b0001110001011011: color_data = 12'b001110100111;
		16'b0001110001011100: color_data = 12'b001110100111;
		16'b0001110001011101: color_data = 12'b001110100111;
		16'b0001110001011110: color_data = 12'b001110100111;
		16'b0001110001011111: color_data = 12'b001110100111;
		16'b0001110001100000: color_data = 12'b001110100111;
		16'b0001110001100001: color_data = 12'b001110100111;
		16'b0001110001100010: color_data = 12'b001110100111;
		16'b0001110001100011: color_data = 12'b001110100111;
		16'b0001110001100100: color_data = 12'b001110100111;
		16'b0001110001100101: color_data = 12'b001110100111;
		16'b0001110001100110: color_data = 12'b001110100111;
		16'b0001110001100111: color_data = 12'b001110100111;
		16'b0001110001101000: color_data = 12'b001110100111;
		16'b0001110001101001: color_data = 12'b001110100111;
		16'b0001110001101010: color_data = 12'b001110100111;
		16'b0001110001101011: color_data = 12'b001110100111;
		16'b0001110001101100: color_data = 12'b001110100111;
		16'b0001110001101101: color_data = 12'b001110100111;
		16'b0001110001101110: color_data = 12'b001110100111;
		16'b0001110001110101: color_data = 12'b001110100111;
		16'b0001110001110110: color_data = 12'b001110100111;
		16'b0001110001110111: color_data = 12'b001110100111;
		16'b0001110001111000: color_data = 12'b001110100111;
		16'b0001110001111001: color_data = 12'b001110100111;
		16'b0001110001111010: color_data = 12'b001110100111;
		16'b0001110001111011: color_data = 12'b001110100111;
		16'b0001110001111100: color_data = 12'b001110100111;
		16'b0001110001111101: color_data = 12'b001110100111;
		16'b0001110001111110: color_data = 12'b001110100111;
		16'b0001110001111111: color_data = 12'b001110100111;
		16'b0001110010000000: color_data = 12'b001110100111;
		16'b0001110010000001: color_data = 12'b001110100111;
		16'b0001110010000010: color_data = 12'b001110100111;
		16'b0001110010000011: color_data = 12'b001110100111;
		16'b0001110010000100: color_data = 12'b001110100111;
		16'b0001110010000101: color_data = 12'b001110100111;
		16'b0001110010000110: color_data = 12'b001110100111;
		16'b0001110010000111: color_data = 12'b001110100111;
		16'b0001110010001000: color_data = 12'b001110100111;
		16'b0001110010001001: color_data = 12'b001110100111;
		16'b0001110010001010: color_data = 12'b001110100111;
		16'b0001110010001011: color_data = 12'b001110100111;
		16'b0001110010001100: color_data = 12'b001110100111;
		16'b0001110010001101: color_data = 12'b001110100111;
		16'b0001110010001110: color_data = 12'b001110100111;
		16'b0001110010001111: color_data = 12'b001110100111;
		16'b0001110010010000: color_data = 12'b001110100111;
		16'b0001110010010001: color_data = 12'b001110100111;
		16'b0001110010010010: color_data = 12'b001110100111;
		16'b0001110010010011: color_data = 12'b001110100111;
		16'b0001110010100110: color_data = 12'b001110100111;
		16'b0001110010100111: color_data = 12'b001110100111;
		16'b0001110010101000: color_data = 12'b001110100111;
		16'b0001110010101001: color_data = 12'b001110100111;
		16'b0001110010101010: color_data = 12'b001110100111;
		16'b0001110010101011: color_data = 12'b001110100111;
		16'b0001110010101100: color_data = 12'b001110100111;
		16'b0001110010101101: color_data = 12'b001110100111;
		16'b0001110010101110: color_data = 12'b001110100111;
		16'b0001110010101111: color_data = 12'b001110100111;
		16'b0001110010110000: color_data = 12'b001110100111;
		16'b0001110010110001: color_data = 12'b001110100111;
		16'b0001110010110010: color_data = 12'b001110100111;
		16'b0001110010110011: color_data = 12'b001110100111;
		16'b0001110010110100: color_data = 12'b001110100111;
		16'b0001110010110101: color_data = 12'b001110100111;
		16'b0001110010110110: color_data = 12'b001110100111;
		16'b0001110010110111: color_data = 12'b001110100111;
		16'b0001110010111000: color_data = 12'b001110100111;
		16'b0001110010111001: color_data = 12'b001110100111;
		16'b0001110010111010: color_data = 12'b001110100111;
		16'b0001110010111011: color_data = 12'b001110100111;
		16'b0001110010111100: color_data = 12'b001110100111;
		16'b0001110010111101: color_data = 12'b001110100111;
		16'b0001110010111110: color_data = 12'b001110100111;
		16'b0001110010111111: color_data = 12'b001110100111;
		16'b0001110011000000: color_data = 12'b001110100111;
		16'b0001110011000001: color_data = 12'b001110100111;
		16'b0001110011000010: color_data = 12'b001110100111;
		16'b0001110011000011: color_data = 12'b001110100111;
		16'b0001110011000100: color_data = 12'b001110100111;
		16'b0001110011001011: color_data = 12'b001110100111;
		16'b0001110011001100: color_data = 12'b001110100111;
		16'b0001110011001101: color_data = 12'b001110100111;
		16'b0001110011001110: color_data = 12'b001110100111;
		16'b0001110011001111: color_data = 12'b001110100111;
		16'b0001110011010000: color_data = 12'b001110100111;
		16'b0001110011010001: color_data = 12'b001110100111;
		16'b0001110011010010: color_data = 12'b001110100111;
		16'b0001110011010011: color_data = 12'b001110100111;
		16'b0001110011010100: color_data = 12'b001110100111;
		16'b0001110011010101: color_data = 12'b001110100111;
		16'b0001110011010110: color_data = 12'b001110100111;
		16'b0001110011010111: color_data = 12'b001110100111;
		16'b0001110011011000: color_data = 12'b001110100111;
		16'b0001110011011001: color_data = 12'b001110100111;
		16'b0001110011011010: color_data = 12'b001110100111;
		16'b0001110011011011: color_data = 12'b001110100111;
		16'b0001110011011100: color_data = 12'b001110100111;
		16'b0001110011011101: color_data = 12'b001110100111;
		16'b0001110011011110: color_data = 12'b001110100111;
		16'b0001110011011111: color_data = 12'b001110100111;
		16'b0001110011100000: color_data = 12'b001110100111;
		16'b0001110011100001: color_data = 12'b001110100111;
		16'b0001110011100010: color_data = 12'b001110100111;
		16'b0001110011100011: color_data = 12'b001110100111;
		16'b0001110011100100: color_data = 12'b001110100111;
		16'b0001110011100101: color_data = 12'b001110100111;
		16'b0001110011100110: color_data = 12'b001110100111;
		16'b0001110011100111: color_data = 12'b001110100111;
		16'b0001110011101000: color_data = 12'b001110100111;
		16'b0001110011101001: color_data = 12'b001110100111;
		16'b0001110011101010: color_data = 12'b001110100111;
		16'b0001110011101011: color_data = 12'b001110100111;
		16'b0001110011101100: color_data = 12'b001110100111;
		16'b0001110011101101: color_data = 12'b001110100111;
		16'b0001110011101110: color_data = 12'b001110100111;
		16'b0001110011101111: color_data = 12'b001110100111;
		16'b0001110011110110: color_data = 12'b001110100111;
		16'b0001110011110111: color_data = 12'b001110100111;
		16'b0001110011111000: color_data = 12'b001110100111;
		16'b0001110011111001: color_data = 12'b001110100111;
		16'b0001110011111010: color_data = 12'b001110100111;
		16'b0001110011111011: color_data = 12'b001110100111;
		16'b0001110011111100: color_data = 12'b001110100111;
		16'b0001110011111101: color_data = 12'b001110100111;
		16'b0001110011111110: color_data = 12'b001110100111;
		16'b0001110011111111: color_data = 12'b001110100111;
		16'b0001110100000000: color_data = 12'b001110100111;
		16'b0001110100000001: color_data = 12'b001110100111;
		16'b0001110100000010: color_data = 12'b001110100111;
		16'b0001110100000011: color_data = 12'b001110100111;
		16'b0001110100000100: color_data = 12'b001110100111;
		16'b0001110100000101: color_data = 12'b001110100111;
		16'b0001110100000110: color_data = 12'b001110100111;
		16'b0001110100000111: color_data = 12'b001110100111;
		16'b0001110100001000: color_data = 12'b001110100111;
		16'b0001110100001001: color_data = 12'b001110100111;
		16'b0001110100001010: color_data = 12'b001110100111;
		16'b0001110100001011: color_data = 12'b001110100111;
		16'b0001110100001100: color_data = 12'b001110100111;
		16'b0001110100001101: color_data = 12'b001110100111;
		16'b0001110100001110: color_data = 12'b001110100111;
		16'b0001110100001111: color_data = 12'b001110100111;
		16'b0001110100010000: color_data = 12'b001110100111;
		16'b0001110100010001: color_data = 12'b001110100111;
		16'b0001110100010010: color_data = 12'b001110100111;
		16'b0001110100010011: color_data = 12'b001110100111;
		16'b0001110100010100: color_data = 12'b001110100111;
		16'b0001110100010101: color_data = 12'b001110100111;
		16'b0001110100010110: color_data = 12'b001110100111;
		16'b0001110100010111: color_data = 12'b001110100111;
		16'b0001110100011000: color_data = 12'b001110100111;
		16'b0001110100011001: color_data = 12'b001110100111;
		16'b0001110100011010: color_data = 12'b001110100111;
		16'b0001110100011011: color_data = 12'b001110100111;
		16'b0001110100011100: color_data = 12'b001110100111;
		16'b0001110100011101: color_data = 12'b001110100111;
		16'b0001110100011110: color_data = 12'b001110100111;
		16'b0001110100011111: color_data = 12'b001110100111;
		16'b0001110100100000: color_data = 12'b001110100111;
		16'b0001110100100001: color_data = 12'b001110100111;
		16'b0001110100100010: color_data = 12'b001110100111;
		16'b0001110100100011: color_data = 12'b001110100111;
		16'b0001110100100100: color_data = 12'b001110100111;
		16'b0001110100100101: color_data = 12'b001110100111;
		16'b0001110100100110: color_data = 12'b001110100111;
		16'b0001110100101101: color_data = 12'b001110100111;
		16'b0001110100101110: color_data = 12'b001110100111;
		16'b0001110100101111: color_data = 12'b001110100111;
		16'b0001110100110000: color_data = 12'b001110100111;
		16'b0001110100110001: color_data = 12'b001110100111;
		16'b0001110100110010: color_data = 12'b001110100111;
		16'b0001110100110011: color_data = 12'b001110100111;
		16'b0001110100110100: color_data = 12'b001110100111;
		16'b0001110100110101: color_data = 12'b001110100111;
		16'b0001110100110110: color_data = 12'b001110100111;
		16'b0001110100110111: color_data = 12'b001110100111;
		16'b0001110100111000: color_data = 12'b001110100111;
		16'b0001110100111001: color_data = 12'b001110100111;
		16'b0001110100111010: color_data = 12'b001110100111;
		16'b0001110100111011: color_data = 12'b001110100111;
		16'b0001110100111100: color_data = 12'b001110100111;
		16'b0001110100111101: color_data = 12'b001110100111;
		16'b0001110100111110: color_data = 12'b001110100111;
		16'b0001110100111111: color_data = 12'b001110100111;
		16'b0001110101000000: color_data = 12'b001110100111;
		16'b0001110101000001: color_data = 12'b001110100111;
		16'b0001110101000010: color_data = 12'b001110100111;
		16'b0001110101000011: color_data = 12'b001110100111;
		16'b0001110101000100: color_data = 12'b001110100111;
		16'b0001110101000101: color_data = 12'b001110100111;
		16'b0001110101000110: color_data = 12'b001110100111;
		16'b0001110101000111: color_data = 12'b001110100111;
		16'b0001110101001000: color_data = 12'b001110100111;
		16'b0001110101001001: color_data = 12'b001110100111;
		16'b0001110101001010: color_data = 12'b001110100111;
		16'b0001110101011110: color_data = 12'b001110100111;
		16'b0001110101011111: color_data = 12'b001110100111;
		16'b0001110101100000: color_data = 12'b001110100111;
		16'b0001110101100001: color_data = 12'b001110100111;
		16'b0001110101100010: color_data = 12'b001110100111;
		16'b0001110101100011: color_data = 12'b001110100111;
		16'b0001110101100100: color_data = 12'b001110100111;
		16'b0001110101100101: color_data = 12'b001110100111;
		16'b0001110101100110: color_data = 12'b001110100111;
		16'b0001110101100111: color_data = 12'b001110100111;
		16'b0001110101101000: color_data = 12'b001110100111;
		16'b0001110101101001: color_data = 12'b001110100111;
		16'b0001110101101010: color_data = 12'b001110100111;
		16'b0001110101101011: color_data = 12'b001110100111;
		16'b0001110101101100: color_data = 12'b001110100111;
		16'b0001110101101101: color_data = 12'b001110100111;
		16'b0001110101101110: color_data = 12'b001110100111;
		16'b0001110101101111: color_data = 12'b001110100111;
		16'b0001110101110000: color_data = 12'b001110100111;
		16'b0001110101110001: color_data = 12'b001110100111;
		16'b0001110101110010: color_data = 12'b001110100111;
		16'b0001110101110011: color_data = 12'b001110100111;
		16'b0001110101110100: color_data = 12'b001110100111;
		16'b0001110101110101: color_data = 12'b001110100111;
		16'b0001110101110110: color_data = 12'b001110100111;
		16'b0001110101110111: color_data = 12'b001110100111;
		16'b0001110101111000: color_data = 12'b001110100111;
		16'b0001110101111001: color_data = 12'b001110100111;
		16'b0001110101111010: color_data = 12'b001110100111;
		16'b0001110101111011: color_data = 12'b001110100111;
		16'b0001111000000111: color_data = 12'b001110100111;
		16'b0001111000001000: color_data = 12'b001110100111;
		16'b0001111000001001: color_data = 12'b001110100111;
		16'b0001111000001010: color_data = 12'b001110100111;
		16'b0001111000001011: color_data = 12'b001110100111;
		16'b0001111000001100: color_data = 12'b001110100111;
		16'b0001111000001101: color_data = 12'b001110100111;
		16'b0001111000001110: color_data = 12'b001110100111;
		16'b0001111000001111: color_data = 12'b001110100111;
		16'b0001111000010000: color_data = 12'b001110100111;
		16'b0001111000010001: color_data = 12'b001110100111;
		16'b0001111000010010: color_data = 12'b001110100111;
		16'b0001111000010011: color_data = 12'b001110100111;
		16'b0001111000010100: color_data = 12'b001110100111;
		16'b0001111000010101: color_data = 12'b001110100111;
		16'b0001111000010110: color_data = 12'b001110100111;
		16'b0001111000010111: color_data = 12'b001110100111;
		16'b0001111000011000: color_data = 12'b001110100111;
		16'b0001111000011001: color_data = 12'b001110100111;
		16'b0001111000011010: color_data = 12'b001110100111;
		16'b0001111000011011: color_data = 12'b001110100111;
		16'b0001111000011100: color_data = 12'b001110100111;
		16'b0001111000011101: color_data = 12'b001110100111;
		16'b0001111000011110: color_data = 12'b001110100111;
		16'b0001111000011111: color_data = 12'b001110100111;
		16'b0001111000100000: color_data = 12'b001110100111;
		16'b0001111000100001: color_data = 12'b001110100111;
		16'b0001111000100010: color_data = 12'b001110100111;
		16'b0001111000100011: color_data = 12'b001110100111;
		16'b0001111000100100: color_data = 12'b001110100111;
		16'b0001111000101011: color_data = 12'b001110100111;
		16'b0001111000101100: color_data = 12'b001110100111;
		16'b0001111000101101: color_data = 12'b001110100111;
		16'b0001111000101110: color_data = 12'b001110100111;
		16'b0001111000101111: color_data = 12'b001110100111;
		16'b0001111000110000: color_data = 12'b001110100111;
		16'b0001111000110001: color_data = 12'b001110100111;
		16'b0001111000110010: color_data = 12'b001110100111;
		16'b0001111000110011: color_data = 12'b001110100111;
		16'b0001111000110100: color_data = 12'b001110100111;
		16'b0001111000110101: color_data = 12'b001110100111;
		16'b0001111000110110: color_data = 12'b001110100111;
		16'b0001111000110111: color_data = 12'b001110100111;
		16'b0001111001000100: color_data = 12'b001110100111;
		16'b0001111001000101: color_data = 12'b001110100111;
		16'b0001111001000110: color_data = 12'b001110100111;
		16'b0001111001000111: color_data = 12'b001110100111;
		16'b0001111001001000: color_data = 12'b001110100111;
		16'b0001111001001001: color_data = 12'b001110100111;
		16'b0001111001001010: color_data = 12'b001110100111;
		16'b0001111001001011: color_data = 12'b001110100111;
		16'b0001111001001100: color_data = 12'b001110100111;
		16'b0001111001001101: color_data = 12'b001110100111;
		16'b0001111001001110: color_data = 12'b001110100111;
		16'b0001111001001111: color_data = 12'b001110100111;
		16'b0001111001010110: color_data = 12'b001110100111;
		16'b0001111001010111: color_data = 12'b001110100111;
		16'b0001111001011000: color_data = 12'b001110100111;
		16'b0001111001011001: color_data = 12'b001110100111;
		16'b0001111001011010: color_data = 12'b001110100111;
		16'b0001111001011011: color_data = 12'b001110100111;
		16'b0001111001011100: color_data = 12'b001110100111;
		16'b0001111001011101: color_data = 12'b001110100111;
		16'b0001111001011110: color_data = 12'b001110100111;
		16'b0001111001011111: color_data = 12'b001110100111;
		16'b0001111001100000: color_data = 12'b001110100111;
		16'b0001111001100001: color_data = 12'b001110100111;
		16'b0001111001100010: color_data = 12'b001110100111;
		16'b0001111001100011: color_data = 12'b001110100111;
		16'b0001111001100100: color_data = 12'b001110100111;
		16'b0001111001100101: color_data = 12'b001110100111;
		16'b0001111001100110: color_data = 12'b001110100111;
		16'b0001111001100111: color_data = 12'b001110100111;
		16'b0001111001101000: color_data = 12'b001110100111;
		16'b0001111001101001: color_data = 12'b001110100111;
		16'b0001111001101010: color_data = 12'b001110100111;
		16'b0001111001101011: color_data = 12'b001110100111;
		16'b0001111001101100: color_data = 12'b001110100111;
		16'b0001111001101101: color_data = 12'b001110100111;
		16'b0001111001101110: color_data = 12'b001110100111;
		16'b0001111001110101: color_data = 12'b001110100111;
		16'b0001111001110110: color_data = 12'b001110100111;
		16'b0001111001110111: color_data = 12'b001110100111;
		16'b0001111001111000: color_data = 12'b001110100111;
		16'b0001111001111001: color_data = 12'b001110100111;
		16'b0001111001111010: color_data = 12'b001110100111;
		16'b0001111001111011: color_data = 12'b001110100111;
		16'b0001111001111100: color_data = 12'b001110100111;
		16'b0001111001111101: color_data = 12'b001110100111;
		16'b0001111001111110: color_data = 12'b001110100111;
		16'b0001111001111111: color_data = 12'b001110100111;
		16'b0001111010000000: color_data = 12'b001110100111;
		16'b0001111010000001: color_data = 12'b001110100111;
		16'b0001111010000010: color_data = 12'b001110100111;
		16'b0001111010000011: color_data = 12'b001110100111;
		16'b0001111010000100: color_data = 12'b001110100111;
		16'b0001111010000101: color_data = 12'b001110100111;
		16'b0001111010000110: color_data = 12'b001110100111;
		16'b0001111010000111: color_data = 12'b001110100111;
		16'b0001111010001000: color_data = 12'b001110100111;
		16'b0001111010001001: color_data = 12'b001110100111;
		16'b0001111010001010: color_data = 12'b001110100111;
		16'b0001111010001011: color_data = 12'b001110100111;
		16'b0001111010001100: color_data = 12'b001110100111;
		16'b0001111010001101: color_data = 12'b001110100111;
		16'b0001111010001110: color_data = 12'b001110100111;
		16'b0001111010001111: color_data = 12'b001110100111;
		16'b0001111010010000: color_data = 12'b001110100111;
		16'b0001111010010001: color_data = 12'b001110100111;
		16'b0001111010010010: color_data = 12'b001110100111;
		16'b0001111010010011: color_data = 12'b001110100111;
		16'b0001111010100110: color_data = 12'b001110100111;
		16'b0001111010100111: color_data = 12'b001110100111;
		16'b0001111010101000: color_data = 12'b001110100111;
		16'b0001111010101001: color_data = 12'b001110100111;
		16'b0001111010101010: color_data = 12'b001110100111;
		16'b0001111010101011: color_data = 12'b001110100111;
		16'b0001111010101100: color_data = 12'b001110100111;
		16'b0001111010101101: color_data = 12'b001110100111;
		16'b0001111010101110: color_data = 12'b001110100111;
		16'b0001111010101111: color_data = 12'b001110100111;
		16'b0001111010110000: color_data = 12'b001110100111;
		16'b0001111010110001: color_data = 12'b001110100111;
		16'b0001111010110010: color_data = 12'b001110100111;
		16'b0001111010110011: color_data = 12'b001110100111;
		16'b0001111010110100: color_data = 12'b001110100111;
		16'b0001111010110101: color_data = 12'b001110100111;
		16'b0001111010110110: color_data = 12'b001110100111;
		16'b0001111010110111: color_data = 12'b001110100111;
		16'b0001111010111000: color_data = 12'b001110100111;
		16'b0001111010111001: color_data = 12'b001110100111;
		16'b0001111010111010: color_data = 12'b001110100111;
		16'b0001111010111011: color_data = 12'b001110100111;
		16'b0001111010111100: color_data = 12'b001110100111;
		16'b0001111010111101: color_data = 12'b001110100111;
		16'b0001111010111110: color_data = 12'b001110100111;
		16'b0001111010111111: color_data = 12'b001110100111;
		16'b0001111011000000: color_data = 12'b001110100111;
		16'b0001111011000001: color_data = 12'b001110100111;
		16'b0001111011000010: color_data = 12'b001110100111;
		16'b0001111011000011: color_data = 12'b001110100111;
		16'b0001111011000100: color_data = 12'b001110100111;
		16'b0001111011001011: color_data = 12'b001110100111;
		16'b0001111011001100: color_data = 12'b001110100111;
		16'b0001111011001101: color_data = 12'b001110100111;
		16'b0001111011001110: color_data = 12'b001110100111;
		16'b0001111011001111: color_data = 12'b001110100111;
		16'b0001111011010000: color_data = 12'b001110100111;
		16'b0001111011010001: color_data = 12'b001110100111;
		16'b0001111011010010: color_data = 12'b001110100111;
		16'b0001111011010011: color_data = 12'b001110100111;
		16'b0001111011010100: color_data = 12'b001110100111;
		16'b0001111011010101: color_data = 12'b001110100111;
		16'b0001111011010110: color_data = 12'b001110100111;
		16'b0001111011010111: color_data = 12'b001110100111;
		16'b0001111011011000: color_data = 12'b001110100111;
		16'b0001111011011001: color_data = 12'b001110100111;
		16'b0001111011011010: color_data = 12'b001110100111;
		16'b0001111011011011: color_data = 12'b001110100111;
		16'b0001111011011100: color_data = 12'b001110100111;
		16'b0001111011011101: color_data = 12'b001110100111;
		16'b0001111011011110: color_data = 12'b001110100111;
		16'b0001111011011111: color_data = 12'b001110100111;
		16'b0001111011100000: color_data = 12'b001110100111;
		16'b0001111011100001: color_data = 12'b001110100111;
		16'b0001111011100010: color_data = 12'b001110100111;
		16'b0001111011100011: color_data = 12'b001110100111;
		16'b0001111011100100: color_data = 12'b001110100111;
		16'b0001111011100101: color_data = 12'b001110100111;
		16'b0001111011100110: color_data = 12'b001110100111;
		16'b0001111011100111: color_data = 12'b001110100111;
		16'b0001111011101000: color_data = 12'b001110100111;
		16'b0001111011101001: color_data = 12'b001110100111;
		16'b0001111011101010: color_data = 12'b001110100111;
		16'b0001111011101011: color_data = 12'b001110100111;
		16'b0001111011101100: color_data = 12'b001110100111;
		16'b0001111011101101: color_data = 12'b001110100111;
		16'b0001111011101110: color_data = 12'b001110100111;
		16'b0001111011101111: color_data = 12'b001110100111;
		16'b0001111011110110: color_data = 12'b001110100111;
		16'b0001111011110111: color_data = 12'b001110100111;
		16'b0001111011111000: color_data = 12'b001110100111;
		16'b0001111011111001: color_data = 12'b001110100111;
		16'b0001111011111010: color_data = 12'b001110100111;
		16'b0001111011111011: color_data = 12'b001110100111;
		16'b0001111011111100: color_data = 12'b001110100111;
		16'b0001111011111101: color_data = 12'b001110100111;
		16'b0001111011111110: color_data = 12'b001110100111;
		16'b0001111011111111: color_data = 12'b001110100111;
		16'b0001111100000000: color_data = 12'b001110100111;
		16'b0001111100000001: color_data = 12'b001110100111;
		16'b0001111100000010: color_data = 12'b001110100111;
		16'b0001111100000011: color_data = 12'b001110100111;
		16'b0001111100000100: color_data = 12'b001110100111;
		16'b0001111100000101: color_data = 12'b001110100111;
		16'b0001111100000110: color_data = 12'b001110100111;
		16'b0001111100000111: color_data = 12'b001110100111;
		16'b0001111100001000: color_data = 12'b001110100111;
		16'b0001111100001001: color_data = 12'b001110100111;
		16'b0001111100001010: color_data = 12'b001110100111;
		16'b0001111100001011: color_data = 12'b001110100111;
		16'b0001111100001100: color_data = 12'b001110100111;
		16'b0001111100001101: color_data = 12'b001110100111;
		16'b0001111100001110: color_data = 12'b001110100111;
		16'b0001111100001111: color_data = 12'b001110100111;
		16'b0001111100010000: color_data = 12'b001110100111;
		16'b0001111100010001: color_data = 12'b001110100111;
		16'b0001111100010010: color_data = 12'b001110100111;
		16'b0001111100010011: color_data = 12'b001110100111;
		16'b0001111100010100: color_data = 12'b001110100111;
		16'b0001111100010101: color_data = 12'b001110100111;
		16'b0001111100010110: color_data = 12'b001110100111;
		16'b0001111100010111: color_data = 12'b001110100111;
		16'b0001111100011000: color_data = 12'b001110100111;
		16'b0001111100011001: color_data = 12'b001110100111;
		16'b0001111100011010: color_data = 12'b001110100111;
		16'b0001111100011011: color_data = 12'b001110100111;
		16'b0001111100011100: color_data = 12'b001110100111;
		16'b0001111100011101: color_data = 12'b001110100111;
		16'b0001111100011110: color_data = 12'b001110100111;
		16'b0001111100011111: color_data = 12'b001110100111;
		16'b0001111100100000: color_data = 12'b001110100111;
		16'b0001111100100001: color_data = 12'b001110100111;
		16'b0001111100100010: color_data = 12'b001110100111;
		16'b0001111100100011: color_data = 12'b001110100111;
		16'b0001111100100100: color_data = 12'b001110100111;
		16'b0001111100100101: color_data = 12'b001110100111;
		16'b0001111100100110: color_data = 12'b001110100111;
		16'b0001111100101101: color_data = 12'b001110100111;
		16'b0001111100101110: color_data = 12'b001110100111;
		16'b0001111100101111: color_data = 12'b001110100111;
		16'b0001111100110000: color_data = 12'b001110100111;
		16'b0001111100110001: color_data = 12'b001110100111;
		16'b0001111100110010: color_data = 12'b001110100111;
		16'b0001111100110011: color_data = 12'b001110100111;
		16'b0001111100110100: color_data = 12'b001110100111;
		16'b0001111100110101: color_data = 12'b001110100111;
		16'b0001111100110110: color_data = 12'b001110100111;
		16'b0001111100110111: color_data = 12'b001110100111;
		16'b0001111100111000: color_data = 12'b001110100111;
		16'b0001111100111001: color_data = 12'b001110100111;
		16'b0001111100111010: color_data = 12'b001110100111;
		16'b0001111100111011: color_data = 12'b001110100111;
		16'b0001111100111100: color_data = 12'b001110100111;
		16'b0001111100111101: color_data = 12'b001110100111;
		16'b0001111100111110: color_data = 12'b001110100111;
		16'b0001111100111111: color_data = 12'b001110100111;
		16'b0001111101000000: color_data = 12'b001110100111;
		16'b0001111101000001: color_data = 12'b001110100111;
		16'b0001111101000010: color_data = 12'b001110100111;
		16'b0001111101000011: color_data = 12'b001110100111;
		16'b0001111101000100: color_data = 12'b001110100111;
		16'b0001111101000101: color_data = 12'b001110100111;
		16'b0001111101000110: color_data = 12'b001110100111;
		16'b0001111101000111: color_data = 12'b001110100111;
		16'b0001111101001000: color_data = 12'b001110100111;
		16'b0001111101001001: color_data = 12'b001110100111;
		16'b0001111101001010: color_data = 12'b001110100111;
		16'b0001111101011110: color_data = 12'b001110100111;
		16'b0001111101011111: color_data = 12'b001110100111;
		16'b0001111101100000: color_data = 12'b001110100111;
		16'b0001111101100001: color_data = 12'b001110100111;
		16'b0001111101100010: color_data = 12'b001110100111;
		16'b0001111101100011: color_data = 12'b001110100111;
		16'b0001111101100100: color_data = 12'b001110100111;
		16'b0001111101100101: color_data = 12'b001110100111;
		16'b0001111101100110: color_data = 12'b001110100111;
		16'b0001111101100111: color_data = 12'b001110100111;
		16'b0001111101101000: color_data = 12'b001110100111;
		16'b0001111101101001: color_data = 12'b001110100111;
		16'b0001111101101010: color_data = 12'b001110100111;
		16'b0001111101101011: color_data = 12'b001110100111;
		16'b0001111101101100: color_data = 12'b001110100111;
		16'b0001111101101101: color_data = 12'b001110100111;
		16'b0001111101101110: color_data = 12'b001110100111;
		16'b0001111101101111: color_data = 12'b001110100111;
		16'b0001111101110000: color_data = 12'b001110100111;
		16'b0001111101110001: color_data = 12'b001110100111;
		16'b0001111101110010: color_data = 12'b001110100111;
		16'b0001111101110011: color_data = 12'b001110100111;
		16'b0001111101110100: color_data = 12'b001110100111;
		16'b0001111101110101: color_data = 12'b001110100111;
		16'b0001111101110110: color_data = 12'b001110100111;
		16'b0001111101110111: color_data = 12'b001110100111;
		16'b0001111101111000: color_data = 12'b001110100111;
		16'b0001111101111001: color_data = 12'b001110100111;
		16'b0001111101111010: color_data = 12'b001110100111;
		16'b0001111101111011: color_data = 12'b001110100111;
		16'b0010000000000111: color_data = 12'b001110100111;
		16'b0010000000001000: color_data = 12'b001110100111;
		16'b0010000000001001: color_data = 12'b001110100111;
		16'b0010000000001010: color_data = 12'b001110100111;
		16'b0010000000001011: color_data = 12'b001110100111;
		16'b0010000000001100: color_data = 12'b001110100111;
		16'b0010000000001101: color_data = 12'b001110100111;
		16'b0010000000001110: color_data = 12'b001110100111;
		16'b0010000000001111: color_data = 12'b001110100111;
		16'b0010000000010000: color_data = 12'b001110100111;
		16'b0010000000010001: color_data = 12'b001110100111;
		16'b0010000000010010: color_data = 12'b001110100111;
		16'b0010000000010011: color_data = 12'b001110100111;
		16'b0010000000010100: color_data = 12'b001110100111;
		16'b0010000000010101: color_data = 12'b001110100111;
		16'b0010000000010110: color_data = 12'b001110100111;
		16'b0010000000010111: color_data = 12'b001110100111;
		16'b0010000000011000: color_data = 12'b001110100111;
		16'b0010000000011001: color_data = 12'b001110100111;
		16'b0010000000011010: color_data = 12'b001110100111;
		16'b0010000000011011: color_data = 12'b001110100111;
		16'b0010000000011100: color_data = 12'b001110100111;
		16'b0010000000011101: color_data = 12'b001110100111;
		16'b0010000000011110: color_data = 12'b001110100111;
		16'b0010000000011111: color_data = 12'b001110100111;
		16'b0010000000100000: color_data = 12'b001110100111;
		16'b0010000000100001: color_data = 12'b001110100111;
		16'b0010000000100010: color_data = 12'b001110100111;
		16'b0010000000100011: color_data = 12'b001110100111;
		16'b0010000000100100: color_data = 12'b001110100111;
		16'b0010000000101011: color_data = 12'b001110100111;
		16'b0010000000101100: color_data = 12'b001110100111;
		16'b0010000000101101: color_data = 12'b001110100111;
		16'b0010000000101110: color_data = 12'b001110100111;
		16'b0010000000101111: color_data = 12'b001110100111;
		16'b0010000000110000: color_data = 12'b001110100111;
		16'b0010000000110001: color_data = 12'b001110100111;
		16'b0010000000110010: color_data = 12'b001110100111;
		16'b0010000000110011: color_data = 12'b001110100111;
		16'b0010000000110100: color_data = 12'b001110100111;
		16'b0010000000110101: color_data = 12'b001110100111;
		16'b0010000000110110: color_data = 12'b001110100111;
		16'b0010000000110111: color_data = 12'b001110100111;
		16'b0010000001000100: color_data = 12'b001110100111;
		16'b0010000001000101: color_data = 12'b001110100111;
		16'b0010000001000110: color_data = 12'b001110100111;
		16'b0010000001000111: color_data = 12'b001110100111;
		16'b0010000001001000: color_data = 12'b001110100111;
		16'b0010000001001001: color_data = 12'b001110100111;
		16'b0010000001001010: color_data = 12'b001110100111;
		16'b0010000001001011: color_data = 12'b001110100111;
		16'b0010000001001100: color_data = 12'b001110100111;
		16'b0010000001001101: color_data = 12'b001110100111;
		16'b0010000001001110: color_data = 12'b001110100111;
		16'b0010000001001111: color_data = 12'b001110100111;
		16'b0010000001010110: color_data = 12'b001110100111;
		16'b0010000001010111: color_data = 12'b001110100111;
		16'b0010000001011000: color_data = 12'b001110100111;
		16'b0010000001011001: color_data = 12'b001110100111;
		16'b0010000001011010: color_data = 12'b001110100111;
		16'b0010000001011011: color_data = 12'b001110100111;
		16'b0010000001011100: color_data = 12'b001110100111;
		16'b0010000001011101: color_data = 12'b001110100111;
		16'b0010000001011110: color_data = 12'b001110100111;
		16'b0010000001011111: color_data = 12'b001110100111;
		16'b0010000001100000: color_data = 12'b001110100111;
		16'b0010000001100001: color_data = 12'b001110100111;
		16'b0010000001100010: color_data = 12'b001110100111;
		16'b0010000001100011: color_data = 12'b001110100111;
		16'b0010000001100100: color_data = 12'b001110100111;
		16'b0010000001100101: color_data = 12'b001110100111;
		16'b0010000001100110: color_data = 12'b001110100111;
		16'b0010000001100111: color_data = 12'b001110100111;
		16'b0010000001101000: color_data = 12'b001110100111;
		16'b0010000001101001: color_data = 12'b001110100111;
		16'b0010000001101010: color_data = 12'b001110100111;
		16'b0010000001101011: color_data = 12'b001110100111;
		16'b0010000001101100: color_data = 12'b001110100111;
		16'b0010000001101101: color_data = 12'b001110100111;
		16'b0010000001101110: color_data = 12'b001110100111;
		16'b0010000001110101: color_data = 12'b001110100111;
		16'b0010000001110110: color_data = 12'b001110100111;
		16'b0010000001110111: color_data = 12'b001110100111;
		16'b0010000001111000: color_data = 12'b001110100111;
		16'b0010000001111001: color_data = 12'b001110100111;
		16'b0010000001111010: color_data = 12'b001110100111;
		16'b0010000001111011: color_data = 12'b001110100111;
		16'b0010000001111100: color_data = 12'b001110100111;
		16'b0010000001111101: color_data = 12'b001110100111;
		16'b0010000001111110: color_data = 12'b001110100111;
		16'b0010000001111111: color_data = 12'b001110100111;
		16'b0010000010000000: color_data = 12'b001110100111;
		16'b0010000010000001: color_data = 12'b001110100111;
		16'b0010000010000010: color_data = 12'b001110100111;
		16'b0010000010000011: color_data = 12'b001110100111;
		16'b0010000010000100: color_data = 12'b001110100111;
		16'b0010000010000101: color_data = 12'b001110100111;
		16'b0010000010000110: color_data = 12'b001110100111;
		16'b0010000010000111: color_data = 12'b001110100111;
		16'b0010000010001000: color_data = 12'b001110100111;
		16'b0010000010001001: color_data = 12'b001110100111;
		16'b0010000010001010: color_data = 12'b001110100111;
		16'b0010000010001011: color_data = 12'b001110100111;
		16'b0010000010001100: color_data = 12'b001110100111;
		16'b0010000010001101: color_data = 12'b001110100111;
		16'b0010000010001110: color_data = 12'b001110100111;
		16'b0010000010001111: color_data = 12'b001110100111;
		16'b0010000010010000: color_data = 12'b001110100111;
		16'b0010000010010001: color_data = 12'b001110100111;
		16'b0010000010010010: color_data = 12'b001110100111;
		16'b0010000010010011: color_data = 12'b001110100111;
		16'b0010000010100110: color_data = 12'b001110100111;
		16'b0010000010100111: color_data = 12'b001110100111;
		16'b0010000010101000: color_data = 12'b001110100111;
		16'b0010000010101001: color_data = 12'b001110100111;
		16'b0010000010101010: color_data = 12'b001110100111;
		16'b0010000010101011: color_data = 12'b001110100111;
		16'b0010000010101100: color_data = 12'b001110100111;
		16'b0010000010101101: color_data = 12'b001110100111;
		16'b0010000010101110: color_data = 12'b001110100111;
		16'b0010000010101111: color_data = 12'b001110100111;
		16'b0010000010110000: color_data = 12'b001110100111;
		16'b0010000010110001: color_data = 12'b001110100111;
		16'b0010000010110010: color_data = 12'b001110100111;
		16'b0010000010110011: color_data = 12'b001110100111;
		16'b0010000010110100: color_data = 12'b001110100111;
		16'b0010000010110101: color_data = 12'b001110100111;
		16'b0010000010110110: color_data = 12'b001110100111;
		16'b0010000010110111: color_data = 12'b001110100111;
		16'b0010000010111000: color_data = 12'b001110100111;
		16'b0010000010111001: color_data = 12'b001110100111;
		16'b0010000010111010: color_data = 12'b001110100111;
		16'b0010000010111011: color_data = 12'b001110100111;
		16'b0010000010111100: color_data = 12'b001110100111;
		16'b0010000010111101: color_data = 12'b001110100111;
		16'b0010000010111110: color_data = 12'b001110100111;
		16'b0010000010111111: color_data = 12'b001110100111;
		16'b0010000011000000: color_data = 12'b001110100111;
		16'b0010000011000001: color_data = 12'b001110100111;
		16'b0010000011000010: color_data = 12'b001110100111;
		16'b0010000011000011: color_data = 12'b001110100111;
		16'b0010000011000100: color_data = 12'b001110100111;
		16'b0010000011001011: color_data = 12'b001110100111;
		16'b0010000011001100: color_data = 12'b001110100111;
		16'b0010000011001101: color_data = 12'b001110100111;
		16'b0010000011001110: color_data = 12'b001110100111;
		16'b0010000011001111: color_data = 12'b001110100111;
		16'b0010000011010000: color_data = 12'b001110100111;
		16'b0010000011010001: color_data = 12'b001110100111;
		16'b0010000011010010: color_data = 12'b001110100111;
		16'b0010000011010011: color_data = 12'b001110100111;
		16'b0010000011010100: color_data = 12'b001110100111;
		16'b0010000011010101: color_data = 12'b001110100111;
		16'b0010000011010110: color_data = 12'b001110100111;
		16'b0010000011010111: color_data = 12'b001110100111;
		16'b0010000011011000: color_data = 12'b001110100111;
		16'b0010000011011001: color_data = 12'b001110100111;
		16'b0010000011011010: color_data = 12'b001110100111;
		16'b0010000011011011: color_data = 12'b001110100111;
		16'b0010000011011100: color_data = 12'b001110100111;
		16'b0010000011011101: color_data = 12'b001110100111;
		16'b0010000011011110: color_data = 12'b001110100111;
		16'b0010000011011111: color_data = 12'b001110100111;
		16'b0010000011100000: color_data = 12'b001110100111;
		16'b0010000011100001: color_data = 12'b001110100111;
		16'b0010000011100010: color_data = 12'b001110100111;
		16'b0010000011100011: color_data = 12'b001110100111;
		16'b0010000011100100: color_data = 12'b001110100111;
		16'b0010000011100101: color_data = 12'b001110100111;
		16'b0010000011100110: color_data = 12'b001110100111;
		16'b0010000011100111: color_data = 12'b001110100111;
		16'b0010000011101000: color_data = 12'b001110100111;
		16'b0010000011101001: color_data = 12'b001110100111;
		16'b0010000011101010: color_data = 12'b001110100111;
		16'b0010000011101011: color_data = 12'b001110100111;
		16'b0010000011101100: color_data = 12'b001110100111;
		16'b0010000011101101: color_data = 12'b001110100111;
		16'b0010000011101110: color_data = 12'b001110100111;
		16'b0010000011101111: color_data = 12'b001110100111;
		16'b0010000011110110: color_data = 12'b001110100111;
		16'b0010000011110111: color_data = 12'b001110100111;
		16'b0010000011111000: color_data = 12'b001110100111;
		16'b0010000011111001: color_data = 12'b001110100111;
		16'b0010000011111010: color_data = 12'b001110100111;
		16'b0010000011111011: color_data = 12'b001110100111;
		16'b0010000011111100: color_data = 12'b001110100111;
		16'b0010000011111101: color_data = 12'b001110100111;
		16'b0010000011111110: color_data = 12'b001110100111;
		16'b0010000011111111: color_data = 12'b001110100111;
		16'b0010000100000000: color_data = 12'b001110100111;
		16'b0010000100000001: color_data = 12'b001110100111;
		16'b0010000100000010: color_data = 12'b001110100111;
		16'b0010000100000011: color_data = 12'b001110100111;
		16'b0010000100000100: color_data = 12'b001110100111;
		16'b0010000100000101: color_data = 12'b001110100111;
		16'b0010000100000110: color_data = 12'b001110100111;
		16'b0010000100000111: color_data = 12'b001110100111;
		16'b0010000100001000: color_data = 12'b001110100111;
		16'b0010000100001001: color_data = 12'b001110100111;
		16'b0010000100001010: color_data = 12'b001110100111;
		16'b0010000100001011: color_data = 12'b001110100111;
		16'b0010000100001100: color_data = 12'b001110100111;
		16'b0010000100001101: color_data = 12'b001110100111;
		16'b0010000100001110: color_data = 12'b001110100111;
		16'b0010000100001111: color_data = 12'b001110100111;
		16'b0010000100010000: color_data = 12'b001110100111;
		16'b0010000100010001: color_data = 12'b001110100111;
		16'b0010000100010010: color_data = 12'b001110100111;
		16'b0010000100010011: color_data = 12'b001110100111;
		16'b0010000100010100: color_data = 12'b001110100111;
		16'b0010000100010101: color_data = 12'b001110100111;
		16'b0010000100010110: color_data = 12'b001110100111;
		16'b0010000100010111: color_data = 12'b001110100111;
		16'b0010000100011000: color_data = 12'b001110100111;
		16'b0010000100011001: color_data = 12'b001110100111;
		16'b0010000100011010: color_data = 12'b001110100111;
		16'b0010000100011011: color_data = 12'b001110100111;
		16'b0010000100011100: color_data = 12'b001110100111;
		16'b0010000100011101: color_data = 12'b001110100111;
		16'b0010000100011110: color_data = 12'b001110100111;
		16'b0010000100011111: color_data = 12'b001110100111;
		16'b0010000100100000: color_data = 12'b001110100111;
		16'b0010000100100001: color_data = 12'b001110100111;
		16'b0010000100100010: color_data = 12'b001110100111;
		16'b0010000100100011: color_data = 12'b001110100111;
		16'b0010000100100100: color_data = 12'b001110100111;
		16'b0010000100100101: color_data = 12'b001110100111;
		16'b0010000100100110: color_data = 12'b001110100111;
		16'b0010000100101101: color_data = 12'b001110100111;
		16'b0010000100101110: color_data = 12'b001110100111;
		16'b0010000100101111: color_data = 12'b001110100111;
		16'b0010000100110000: color_data = 12'b001110100111;
		16'b0010000100110001: color_data = 12'b001110100111;
		16'b0010000100110010: color_data = 12'b001110100111;
		16'b0010000100110011: color_data = 12'b001110100111;
		16'b0010000100110100: color_data = 12'b001110100111;
		16'b0010000100110101: color_data = 12'b001110100111;
		16'b0010000100110110: color_data = 12'b001110100111;
		16'b0010000100110111: color_data = 12'b001110100111;
		16'b0010000100111000: color_data = 12'b001110100111;
		16'b0010000100111001: color_data = 12'b001110100111;
		16'b0010000100111010: color_data = 12'b001110100111;
		16'b0010000100111011: color_data = 12'b001110100111;
		16'b0010000100111100: color_data = 12'b001110100111;
		16'b0010000100111101: color_data = 12'b001110100111;
		16'b0010000100111110: color_data = 12'b001110100111;
		16'b0010000100111111: color_data = 12'b001110100111;
		16'b0010000101000000: color_data = 12'b001110100111;
		16'b0010000101000001: color_data = 12'b001110100111;
		16'b0010000101000010: color_data = 12'b001110100111;
		16'b0010000101000011: color_data = 12'b001110100111;
		16'b0010000101000100: color_data = 12'b001110100111;
		16'b0010000101000101: color_data = 12'b001110100111;
		16'b0010000101000110: color_data = 12'b001110100111;
		16'b0010000101000111: color_data = 12'b001110100111;
		16'b0010000101001000: color_data = 12'b001110100111;
		16'b0010000101001001: color_data = 12'b001110100111;
		16'b0010000101001010: color_data = 12'b001110100111;
		16'b0010000101011110: color_data = 12'b001110100111;
		16'b0010000101011111: color_data = 12'b001110100111;
		16'b0010000101100000: color_data = 12'b001110100111;
		16'b0010000101100001: color_data = 12'b001110100111;
		16'b0010000101100010: color_data = 12'b001110100111;
		16'b0010000101100011: color_data = 12'b001110100111;
		16'b0010000101100100: color_data = 12'b001110100111;
		16'b0010000101100101: color_data = 12'b001110100111;
		16'b0010000101100110: color_data = 12'b001110100111;
		16'b0010000101100111: color_data = 12'b001110100111;
		16'b0010000101101000: color_data = 12'b001110100111;
		16'b0010000101101001: color_data = 12'b001110100111;
		16'b0010000101101010: color_data = 12'b001110100111;
		16'b0010000101101011: color_data = 12'b001110100111;
		16'b0010000101101100: color_data = 12'b001110100111;
		16'b0010000101101101: color_data = 12'b001110100111;
		16'b0010000101101110: color_data = 12'b001110100111;
		16'b0010000101101111: color_data = 12'b001110100111;
		16'b0010000101110000: color_data = 12'b001110100111;
		16'b0010000101110001: color_data = 12'b001110100111;
		16'b0010000101110010: color_data = 12'b001110100111;
		16'b0010000101110011: color_data = 12'b001110100111;
		16'b0010000101110100: color_data = 12'b001110100111;
		16'b0010000101110101: color_data = 12'b001110100111;
		16'b0010000101110110: color_data = 12'b001110100111;
		16'b0010000101110111: color_data = 12'b001110100111;
		16'b0010000101111000: color_data = 12'b001110100111;
		16'b0010000101111001: color_data = 12'b001110100111;
		16'b0010000101111010: color_data = 12'b001110100111;
		16'b0010000101111011: color_data = 12'b001110100111;
		16'b0010001000000111: color_data = 12'b001110100111;
		16'b0010001000001000: color_data = 12'b001110100111;
		16'b0010001000001001: color_data = 12'b001110100111;
		16'b0010001000001010: color_data = 12'b001110100111;
		16'b0010001000001011: color_data = 12'b001110100111;
		16'b0010001000001100: color_data = 12'b001110100111;
		16'b0010001000001101: color_data = 12'b001110100111;
		16'b0010001000001110: color_data = 12'b001110100111;
		16'b0010001000001111: color_data = 12'b001110100111;
		16'b0010001000010000: color_data = 12'b001110100111;
		16'b0010001000010001: color_data = 12'b001110100111;
		16'b0010001000010010: color_data = 12'b001110100111;
		16'b0010001000010011: color_data = 12'b001110100111;
		16'b0010001000010100: color_data = 12'b001110100111;
		16'b0010001000010101: color_data = 12'b001110100111;
		16'b0010001000010110: color_data = 12'b001110100111;
		16'b0010001000010111: color_data = 12'b001110100111;
		16'b0010001000011000: color_data = 12'b001110100111;
		16'b0010001000011001: color_data = 12'b001110100111;
		16'b0010001000011010: color_data = 12'b001110100111;
		16'b0010001000011011: color_data = 12'b001110100111;
		16'b0010001000011100: color_data = 12'b001110100111;
		16'b0010001000011101: color_data = 12'b001110100111;
		16'b0010001000011110: color_data = 12'b001110100111;
		16'b0010001000011111: color_data = 12'b001110100111;
		16'b0010001000100000: color_data = 12'b001110100111;
		16'b0010001000100001: color_data = 12'b001110100111;
		16'b0010001000100010: color_data = 12'b001110100111;
		16'b0010001000100011: color_data = 12'b001110100111;
		16'b0010001000100100: color_data = 12'b001110100111;
		16'b0010001000101011: color_data = 12'b001110100111;
		16'b0010001000101100: color_data = 12'b001110100111;
		16'b0010001000101101: color_data = 12'b001110100111;
		16'b0010001000101110: color_data = 12'b001110100111;
		16'b0010001000101111: color_data = 12'b001110100111;
		16'b0010001000110000: color_data = 12'b001110100111;
		16'b0010001000110001: color_data = 12'b001110100111;
		16'b0010001000110010: color_data = 12'b001110100111;
		16'b0010001000110011: color_data = 12'b001110100111;
		16'b0010001000110100: color_data = 12'b001110100111;
		16'b0010001000110101: color_data = 12'b001110100111;
		16'b0010001000110110: color_data = 12'b001110100111;
		16'b0010001000110111: color_data = 12'b001110100111;
		16'b0010001001000100: color_data = 12'b001110100111;
		16'b0010001001000101: color_data = 12'b001110100111;
		16'b0010001001000110: color_data = 12'b001110100111;
		16'b0010001001000111: color_data = 12'b001110100111;
		16'b0010001001001000: color_data = 12'b001110100111;
		16'b0010001001001001: color_data = 12'b001110100111;
		16'b0010001001001010: color_data = 12'b001110100111;
		16'b0010001001001011: color_data = 12'b001110100111;
		16'b0010001001001100: color_data = 12'b001110100111;
		16'b0010001001001101: color_data = 12'b001110100111;
		16'b0010001001001110: color_data = 12'b001110100111;
		16'b0010001001001111: color_data = 12'b001110100111;
		16'b0010001001010110: color_data = 12'b001110100111;
		16'b0010001001010111: color_data = 12'b001110100111;
		16'b0010001001011000: color_data = 12'b001110100111;
		16'b0010001001011001: color_data = 12'b001110100111;
		16'b0010001001011010: color_data = 12'b001110100111;
		16'b0010001001011011: color_data = 12'b001110100111;
		16'b0010001001011100: color_data = 12'b001110100111;
		16'b0010001001011101: color_data = 12'b001110100111;
		16'b0010001001011110: color_data = 12'b001110100111;
		16'b0010001001011111: color_data = 12'b001110100111;
		16'b0010001001100000: color_data = 12'b001110100111;
		16'b0010001001100001: color_data = 12'b001110100111;
		16'b0010001001100010: color_data = 12'b001110100111;
		16'b0010001001100011: color_data = 12'b001110100111;
		16'b0010001001100100: color_data = 12'b001110100111;
		16'b0010001001100101: color_data = 12'b001110100111;
		16'b0010001001100110: color_data = 12'b001110100111;
		16'b0010001001100111: color_data = 12'b001110100111;
		16'b0010001001101000: color_data = 12'b001110100111;
		16'b0010001001101001: color_data = 12'b001110100111;
		16'b0010001001101010: color_data = 12'b001110100111;
		16'b0010001001101011: color_data = 12'b001110100111;
		16'b0010001001101100: color_data = 12'b001110100111;
		16'b0010001001101101: color_data = 12'b001110100111;
		16'b0010001001101110: color_data = 12'b001110100111;
		16'b0010001001110101: color_data = 12'b001110100111;
		16'b0010001001110110: color_data = 12'b001110100111;
		16'b0010001001110111: color_data = 12'b001110100111;
		16'b0010001001111000: color_data = 12'b001110100111;
		16'b0010001001111001: color_data = 12'b001110100111;
		16'b0010001001111010: color_data = 12'b001110100111;
		16'b0010001001111011: color_data = 12'b001110100111;
		16'b0010001001111100: color_data = 12'b001110100111;
		16'b0010001001111101: color_data = 12'b001110100111;
		16'b0010001001111110: color_data = 12'b001110100111;
		16'b0010001001111111: color_data = 12'b001110100111;
		16'b0010001010000000: color_data = 12'b001110100111;
		16'b0010001010000001: color_data = 12'b001110100111;
		16'b0010001010000010: color_data = 12'b001110100111;
		16'b0010001010000011: color_data = 12'b001110100111;
		16'b0010001010000100: color_data = 12'b001110100111;
		16'b0010001010000101: color_data = 12'b001110100111;
		16'b0010001010000110: color_data = 12'b001110100111;
		16'b0010001010000111: color_data = 12'b001110100111;
		16'b0010001010001000: color_data = 12'b001110100111;
		16'b0010001010001001: color_data = 12'b001110100111;
		16'b0010001010001010: color_data = 12'b001110100111;
		16'b0010001010001011: color_data = 12'b001110100111;
		16'b0010001010001100: color_data = 12'b001110100111;
		16'b0010001010001101: color_data = 12'b001110100111;
		16'b0010001010001110: color_data = 12'b001110100111;
		16'b0010001010001111: color_data = 12'b001110100111;
		16'b0010001010010000: color_data = 12'b001110100111;
		16'b0010001010010001: color_data = 12'b001110100111;
		16'b0010001010010010: color_data = 12'b001110100111;
		16'b0010001010010011: color_data = 12'b001110100111;
		16'b0010001010100110: color_data = 12'b001110100111;
		16'b0010001010100111: color_data = 12'b001110100111;
		16'b0010001010101000: color_data = 12'b001110100111;
		16'b0010001010101001: color_data = 12'b001110100111;
		16'b0010001010101010: color_data = 12'b001110100111;
		16'b0010001010101011: color_data = 12'b001110100111;
		16'b0010001010101100: color_data = 12'b001110100111;
		16'b0010001010101101: color_data = 12'b001110100111;
		16'b0010001010101110: color_data = 12'b001110100111;
		16'b0010001010101111: color_data = 12'b001110100111;
		16'b0010001010110000: color_data = 12'b001110100111;
		16'b0010001010110001: color_data = 12'b001110100111;
		16'b0010001010110010: color_data = 12'b001110100111;
		16'b0010001010110011: color_data = 12'b001110100111;
		16'b0010001010110100: color_data = 12'b001110100111;
		16'b0010001010110101: color_data = 12'b001110100111;
		16'b0010001010110110: color_data = 12'b001110100111;
		16'b0010001010110111: color_data = 12'b001110100111;
		16'b0010001010111000: color_data = 12'b001110100111;
		16'b0010001010111001: color_data = 12'b001110100111;
		16'b0010001010111010: color_data = 12'b001110100111;
		16'b0010001010111011: color_data = 12'b001110100111;
		16'b0010001010111100: color_data = 12'b001110100111;
		16'b0010001010111101: color_data = 12'b001110100111;
		16'b0010001010111110: color_data = 12'b001110100111;
		16'b0010001010111111: color_data = 12'b001110100111;
		16'b0010001011000000: color_data = 12'b001110100111;
		16'b0010001011000001: color_data = 12'b001110100111;
		16'b0010001011000010: color_data = 12'b001110100111;
		16'b0010001011000011: color_data = 12'b001110100111;
		16'b0010001011000100: color_data = 12'b001110100111;
		16'b0010001011001011: color_data = 12'b001110100111;
		16'b0010001011001100: color_data = 12'b001110100111;
		16'b0010001011001101: color_data = 12'b001110100111;
		16'b0010001011001110: color_data = 12'b001110100111;
		16'b0010001011001111: color_data = 12'b001110100111;
		16'b0010001011010000: color_data = 12'b001110100111;
		16'b0010001011010001: color_data = 12'b001110100111;
		16'b0010001011010010: color_data = 12'b001110100111;
		16'b0010001011010011: color_data = 12'b001110100111;
		16'b0010001011010100: color_data = 12'b001110100111;
		16'b0010001011010101: color_data = 12'b001110100111;
		16'b0010001011010110: color_data = 12'b001110100111;
		16'b0010001011010111: color_data = 12'b001110100111;
		16'b0010001011011000: color_data = 12'b001110100111;
		16'b0010001011011001: color_data = 12'b001110100111;
		16'b0010001011011010: color_data = 12'b001110100111;
		16'b0010001011011011: color_data = 12'b001110100111;
		16'b0010001011011100: color_data = 12'b001110100111;
		16'b0010001011011101: color_data = 12'b001110100111;
		16'b0010001011011110: color_data = 12'b001110100111;
		16'b0010001011011111: color_data = 12'b001110100111;
		16'b0010001011100000: color_data = 12'b001110100111;
		16'b0010001011100001: color_data = 12'b001110100111;
		16'b0010001011100010: color_data = 12'b001110100111;
		16'b0010001011100011: color_data = 12'b001110100111;
		16'b0010001011100100: color_data = 12'b001110100111;
		16'b0010001011100101: color_data = 12'b001110100111;
		16'b0010001011100110: color_data = 12'b001110100111;
		16'b0010001011100111: color_data = 12'b001110100111;
		16'b0010001011101000: color_data = 12'b001110100111;
		16'b0010001011101001: color_data = 12'b001110100111;
		16'b0010001011101010: color_data = 12'b001110100111;
		16'b0010001011101011: color_data = 12'b001110100111;
		16'b0010001011101100: color_data = 12'b001110100111;
		16'b0010001011101101: color_data = 12'b001110100111;
		16'b0010001011101110: color_data = 12'b001110100111;
		16'b0010001011101111: color_data = 12'b001110100111;
		16'b0010001011110110: color_data = 12'b001110100111;
		16'b0010001011110111: color_data = 12'b001110100111;
		16'b0010001011111000: color_data = 12'b001110100111;
		16'b0010001011111001: color_data = 12'b001110100111;
		16'b0010001011111010: color_data = 12'b001110100111;
		16'b0010001011111011: color_data = 12'b001110100111;
		16'b0010001011111100: color_data = 12'b001110100111;
		16'b0010001011111101: color_data = 12'b001110100111;
		16'b0010001011111110: color_data = 12'b001110100111;
		16'b0010001011111111: color_data = 12'b001110100111;
		16'b0010001100000000: color_data = 12'b001110100111;
		16'b0010001100000001: color_data = 12'b001110100111;
		16'b0010001100000010: color_data = 12'b001110100111;
		16'b0010001100000011: color_data = 12'b001110100111;
		16'b0010001100000100: color_data = 12'b001110100111;
		16'b0010001100000101: color_data = 12'b001110100111;
		16'b0010001100000110: color_data = 12'b001110100111;
		16'b0010001100000111: color_data = 12'b001110100111;
		16'b0010001100001000: color_data = 12'b001110100111;
		16'b0010001100001001: color_data = 12'b001110100111;
		16'b0010001100001010: color_data = 12'b001110100111;
		16'b0010001100001011: color_data = 12'b001110100111;
		16'b0010001100001100: color_data = 12'b001110100111;
		16'b0010001100001101: color_data = 12'b001110100111;
		16'b0010001100001110: color_data = 12'b001110100111;
		16'b0010001100001111: color_data = 12'b001110100111;
		16'b0010001100010000: color_data = 12'b001110100111;
		16'b0010001100010001: color_data = 12'b001110100111;
		16'b0010001100010010: color_data = 12'b001110100111;
		16'b0010001100010011: color_data = 12'b001110100111;
		16'b0010001100010100: color_data = 12'b001110100111;
		16'b0010001100010101: color_data = 12'b001110100111;
		16'b0010001100010110: color_data = 12'b001110100111;
		16'b0010001100010111: color_data = 12'b001110100111;
		16'b0010001100011000: color_data = 12'b001110100111;
		16'b0010001100011001: color_data = 12'b001110100111;
		16'b0010001100011010: color_data = 12'b001110100111;
		16'b0010001100011011: color_data = 12'b001110100111;
		16'b0010001100011100: color_data = 12'b001110100111;
		16'b0010001100011101: color_data = 12'b001110100111;
		16'b0010001100011110: color_data = 12'b001110100111;
		16'b0010001100011111: color_data = 12'b001110100111;
		16'b0010001100100000: color_data = 12'b001110100111;
		16'b0010001100100001: color_data = 12'b001110100111;
		16'b0010001100100010: color_data = 12'b001110100111;
		16'b0010001100100011: color_data = 12'b001110100111;
		16'b0010001100100100: color_data = 12'b001110100111;
		16'b0010001100100101: color_data = 12'b001110100111;
		16'b0010001100100110: color_data = 12'b001110100111;
		16'b0010001100101101: color_data = 12'b001110100111;
		16'b0010001100101110: color_data = 12'b001110100111;
		16'b0010001100101111: color_data = 12'b001110100111;
		16'b0010001100110000: color_data = 12'b001110100111;
		16'b0010001100110001: color_data = 12'b001110100111;
		16'b0010001100110010: color_data = 12'b001110100111;
		16'b0010001100110011: color_data = 12'b001110100111;
		16'b0010001100110100: color_data = 12'b001110100111;
		16'b0010001100110101: color_data = 12'b001110100111;
		16'b0010001100110110: color_data = 12'b001110100111;
		16'b0010001100110111: color_data = 12'b001110100111;
		16'b0010001100111000: color_data = 12'b001110100111;
		16'b0010001100111001: color_data = 12'b001110100111;
		16'b0010001100111010: color_data = 12'b001110100111;
		16'b0010001100111011: color_data = 12'b001110100111;
		16'b0010001100111100: color_data = 12'b001110100111;
		16'b0010001100111101: color_data = 12'b001110100111;
		16'b0010001100111110: color_data = 12'b001110100111;
		16'b0010001100111111: color_data = 12'b001110100111;
		16'b0010001101000000: color_data = 12'b001110100111;
		16'b0010001101000001: color_data = 12'b001110100111;
		16'b0010001101000010: color_data = 12'b001110100111;
		16'b0010001101000011: color_data = 12'b001110100111;
		16'b0010001101000100: color_data = 12'b001110100111;
		16'b0010001101000101: color_data = 12'b001110100111;
		16'b0010001101000110: color_data = 12'b001110100111;
		16'b0010001101000111: color_data = 12'b001110100111;
		16'b0010001101001000: color_data = 12'b001110100111;
		16'b0010001101001001: color_data = 12'b001110100111;
		16'b0010001101001010: color_data = 12'b001110100111;
		16'b0010001101011110: color_data = 12'b001110100111;
		16'b0010001101011111: color_data = 12'b001110100111;
		16'b0010001101100000: color_data = 12'b001110100111;
		16'b0010001101100001: color_data = 12'b001110100111;
		16'b0010001101100010: color_data = 12'b001110100111;
		16'b0010001101100011: color_data = 12'b001110100111;
		16'b0010001101100100: color_data = 12'b001110100111;
		16'b0010001101100101: color_data = 12'b001110100111;
		16'b0010001101100110: color_data = 12'b001110100111;
		16'b0010001101100111: color_data = 12'b001110100111;
		16'b0010001101101000: color_data = 12'b001110100111;
		16'b0010001101101001: color_data = 12'b001110100111;
		16'b0010001101101010: color_data = 12'b001110100111;
		16'b0010001101101011: color_data = 12'b001110100111;
		16'b0010001101101100: color_data = 12'b001110100111;
		16'b0010001101101101: color_data = 12'b001110100111;
		16'b0010001101101110: color_data = 12'b001110100111;
		16'b0010001101101111: color_data = 12'b001110100111;
		16'b0010001101110000: color_data = 12'b001110100111;
		16'b0010001101110001: color_data = 12'b001110100111;
		16'b0010001101110010: color_data = 12'b001110100111;
		16'b0010001101110011: color_data = 12'b001110100111;
		16'b0010001101110100: color_data = 12'b001110100111;
		16'b0010001101110101: color_data = 12'b001110100111;
		16'b0010001101110110: color_data = 12'b001110100111;
		16'b0010001101110111: color_data = 12'b001110100111;
		16'b0010001101111000: color_data = 12'b001110100111;
		16'b0010001101111001: color_data = 12'b001110100111;
		16'b0010001101111010: color_data = 12'b001110100111;
		16'b0010001101111011: color_data = 12'b001110100111;
		16'b0010010000000111: color_data = 12'b001110100111;
		16'b0010010000001000: color_data = 12'b001110100111;
		16'b0010010000001001: color_data = 12'b001110100111;
		16'b0010010000001010: color_data = 12'b001110100111;
		16'b0010010000001011: color_data = 12'b001110100111;
		16'b0010010000001100: color_data = 12'b001110100111;
		16'b0010010000001101: color_data = 12'b001110100111;
		16'b0010010000001110: color_data = 12'b001110100111;
		16'b0010010000001111: color_data = 12'b001110100111;
		16'b0010010000010000: color_data = 12'b001110100111;
		16'b0010010000010001: color_data = 12'b001110100111;
		16'b0010010000010010: color_data = 12'b001110100111;
		16'b0010010000010011: color_data = 12'b001110100111;
		16'b0010010000010100: color_data = 12'b001110100111;
		16'b0010010000010101: color_data = 12'b001110100111;
		16'b0010010000010110: color_data = 12'b001110100111;
		16'b0010010000010111: color_data = 12'b001110100111;
		16'b0010010000011000: color_data = 12'b001110100111;
		16'b0010010000011001: color_data = 12'b001110100111;
		16'b0010010000011010: color_data = 12'b001110100111;
		16'b0010010000011011: color_data = 12'b001110100111;
		16'b0010010000011100: color_data = 12'b001110100111;
		16'b0010010000011101: color_data = 12'b001110100111;
		16'b0010010000011110: color_data = 12'b001110100111;
		16'b0010010000011111: color_data = 12'b001110100111;
		16'b0010010000100000: color_data = 12'b001110100111;
		16'b0010010000100001: color_data = 12'b001110100111;
		16'b0010010000100010: color_data = 12'b001110100111;
		16'b0010010000100011: color_data = 12'b001110100111;
		16'b0010010000100100: color_data = 12'b001110100111;
		16'b0010010000101011: color_data = 12'b001110100111;
		16'b0010010000101100: color_data = 12'b001110100111;
		16'b0010010000101101: color_data = 12'b001110100111;
		16'b0010010000101110: color_data = 12'b001110100111;
		16'b0010010000101111: color_data = 12'b001110100111;
		16'b0010010000110000: color_data = 12'b001110100111;
		16'b0010010000110001: color_data = 12'b001110100111;
		16'b0010010000110010: color_data = 12'b001110100111;
		16'b0010010000110011: color_data = 12'b001110100111;
		16'b0010010000110100: color_data = 12'b001110100111;
		16'b0010010000110101: color_data = 12'b001110100111;
		16'b0010010000110110: color_data = 12'b001110100111;
		16'b0010010000110111: color_data = 12'b001110100111;
		16'b0010010001000100: color_data = 12'b001110100111;
		16'b0010010001000101: color_data = 12'b001110100111;
		16'b0010010001000110: color_data = 12'b001110100111;
		16'b0010010001000111: color_data = 12'b001110100111;
		16'b0010010001001000: color_data = 12'b001110100111;
		16'b0010010001001001: color_data = 12'b001110100111;
		16'b0010010001001010: color_data = 12'b001110100111;
		16'b0010010001001011: color_data = 12'b001110100111;
		16'b0010010001001100: color_data = 12'b001110100111;
		16'b0010010001001101: color_data = 12'b001110100111;
		16'b0010010001001110: color_data = 12'b001110100111;
		16'b0010010001001111: color_data = 12'b001110100111;
		16'b0010010001010110: color_data = 12'b001110100111;
		16'b0010010001010111: color_data = 12'b001110100111;
		16'b0010010001011000: color_data = 12'b001110100111;
		16'b0010010001011001: color_data = 12'b001110100111;
		16'b0010010001011010: color_data = 12'b001110100111;
		16'b0010010001011011: color_data = 12'b001110100111;
		16'b0010010001011100: color_data = 12'b001110100111;
		16'b0010010001011101: color_data = 12'b001110100111;
		16'b0010010001011110: color_data = 12'b001110100111;
		16'b0010010001011111: color_data = 12'b001110100111;
		16'b0010010001100000: color_data = 12'b001110100111;
		16'b0010010001100001: color_data = 12'b001110100111;
		16'b0010010001100010: color_data = 12'b001110100111;
		16'b0010010001100011: color_data = 12'b001110100111;
		16'b0010010001100100: color_data = 12'b001110100111;
		16'b0010010001100101: color_data = 12'b001110100111;
		16'b0010010001100110: color_data = 12'b001110100111;
		16'b0010010001100111: color_data = 12'b001110100111;
		16'b0010010001101000: color_data = 12'b001110100111;
		16'b0010010001101001: color_data = 12'b001110100111;
		16'b0010010001101010: color_data = 12'b001110100111;
		16'b0010010001101011: color_data = 12'b001110100111;
		16'b0010010001101100: color_data = 12'b001110100111;
		16'b0010010001101101: color_data = 12'b001110100111;
		16'b0010010001101110: color_data = 12'b001110100111;
		16'b0010010001110101: color_data = 12'b001110100111;
		16'b0010010001110110: color_data = 12'b001110100111;
		16'b0010010001110111: color_data = 12'b001110100111;
		16'b0010010001111000: color_data = 12'b001110100111;
		16'b0010010001111001: color_data = 12'b001110100111;
		16'b0010010001111010: color_data = 12'b001110100111;
		16'b0010010001111011: color_data = 12'b001110100111;
		16'b0010010001111100: color_data = 12'b001110100111;
		16'b0010010001111101: color_data = 12'b001110100111;
		16'b0010010001111110: color_data = 12'b001110100111;
		16'b0010010001111111: color_data = 12'b001110100111;
		16'b0010010010000000: color_data = 12'b001110100111;
		16'b0010010010000001: color_data = 12'b001110100111;
		16'b0010010010000010: color_data = 12'b001110100111;
		16'b0010010010000011: color_data = 12'b001110100111;
		16'b0010010010000100: color_data = 12'b001110100111;
		16'b0010010010000101: color_data = 12'b001110100111;
		16'b0010010010000110: color_data = 12'b001110100111;
		16'b0010010010000111: color_data = 12'b001110100111;
		16'b0010010010001000: color_data = 12'b001110100111;
		16'b0010010010001001: color_data = 12'b001110100111;
		16'b0010010010001010: color_data = 12'b001110100111;
		16'b0010010010001011: color_data = 12'b001110100111;
		16'b0010010010001100: color_data = 12'b001110100111;
		16'b0010010010001101: color_data = 12'b001110100111;
		16'b0010010010001110: color_data = 12'b001110100111;
		16'b0010010010001111: color_data = 12'b001110100111;
		16'b0010010010010000: color_data = 12'b001110100111;
		16'b0010010010010001: color_data = 12'b001110100111;
		16'b0010010010010010: color_data = 12'b001110100111;
		16'b0010010010010011: color_data = 12'b001110100111;
		16'b0010010010100110: color_data = 12'b001110100111;
		16'b0010010010100111: color_data = 12'b001110100111;
		16'b0010010010101000: color_data = 12'b001110100111;
		16'b0010010010101001: color_data = 12'b001110100111;
		16'b0010010010101010: color_data = 12'b001110100111;
		16'b0010010010101011: color_data = 12'b001110100111;
		16'b0010010010101100: color_data = 12'b001110100111;
		16'b0010010010101101: color_data = 12'b001110100111;
		16'b0010010010101110: color_data = 12'b001110100111;
		16'b0010010010101111: color_data = 12'b001110100111;
		16'b0010010010110000: color_data = 12'b001110100111;
		16'b0010010010110001: color_data = 12'b001110100111;
		16'b0010010010110010: color_data = 12'b001110100111;
		16'b0010010010110011: color_data = 12'b001110100111;
		16'b0010010010110100: color_data = 12'b001110100111;
		16'b0010010010110101: color_data = 12'b001110100111;
		16'b0010010010110110: color_data = 12'b001110100111;
		16'b0010010010110111: color_data = 12'b001110100111;
		16'b0010010010111000: color_data = 12'b001110100111;
		16'b0010010010111001: color_data = 12'b001110100111;
		16'b0010010010111010: color_data = 12'b001110100111;
		16'b0010010010111011: color_data = 12'b001110100111;
		16'b0010010010111100: color_data = 12'b001110100111;
		16'b0010010010111101: color_data = 12'b001110100111;
		16'b0010010010111110: color_data = 12'b001110100111;
		16'b0010010010111111: color_data = 12'b001110100111;
		16'b0010010011000000: color_data = 12'b001110100111;
		16'b0010010011000001: color_data = 12'b001110100111;
		16'b0010010011000010: color_data = 12'b001110100111;
		16'b0010010011000011: color_data = 12'b001110100111;
		16'b0010010011000100: color_data = 12'b001110100111;
		16'b0010010011001011: color_data = 12'b001110100111;
		16'b0010010011001100: color_data = 12'b001110100111;
		16'b0010010011001101: color_data = 12'b001110100111;
		16'b0010010011001110: color_data = 12'b001110100111;
		16'b0010010011001111: color_data = 12'b001110100111;
		16'b0010010011010000: color_data = 12'b001110100111;
		16'b0010010011010001: color_data = 12'b001110100111;
		16'b0010010011010010: color_data = 12'b001110100111;
		16'b0010010011010011: color_data = 12'b001110100111;
		16'b0010010011010100: color_data = 12'b001110100111;
		16'b0010010011010101: color_data = 12'b001110100111;
		16'b0010010011010110: color_data = 12'b001110100111;
		16'b0010010011010111: color_data = 12'b001110100111;
		16'b0010010011011000: color_data = 12'b001110100111;
		16'b0010010011011001: color_data = 12'b001110100111;
		16'b0010010011011010: color_data = 12'b001110100111;
		16'b0010010011011011: color_data = 12'b001110100111;
		16'b0010010011011100: color_data = 12'b001110100111;
		16'b0010010011011101: color_data = 12'b001110100111;
		16'b0010010011011110: color_data = 12'b001110100111;
		16'b0010010011011111: color_data = 12'b001110100111;
		16'b0010010011100000: color_data = 12'b001110100111;
		16'b0010010011100001: color_data = 12'b001110100111;
		16'b0010010011100010: color_data = 12'b001110100111;
		16'b0010010011100011: color_data = 12'b001110100111;
		16'b0010010011100100: color_data = 12'b001110100111;
		16'b0010010011100101: color_data = 12'b001110100111;
		16'b0010010011100110: color_data = 12'b001110100111;
		16'b0010010011100111: color_data = 12'b001110100111;
		16'b0010010011101000: color_data = 12'b001110100111;
		16'b0010010011101001: color_data = 12'b001110100111;
		16'b0010010011101010: color_data = 12'b001110100111;
		16'b0010010011101011: color_data = 12'b001110100111;
		16'b0010010011101100: color_data = 12'b001110100111;
		16'b0010010011101101: color_data = 12'b001110100111;
		16'b0010010011101110: color_data = 12'b001110100111;
		16'b0010010011101111: color_data = 12'b001110100111;
		16'b0010010011110110: color_data = 12'b001110100111;
		16'b0010010011110111: color_data = 12'b001110100111;
		16'b0010010011111000: color_data = 12'b001110100111;
		16'b0010010011111001: color_data = 12'b001110100111;
		16'b0010010011111010: color_data = 12'b001110100111;
		16'b0010010011111011: color_data = 12'b001110100111;
		16'b0010010011111100: color_data = 12'b001110100111;
		16'b0010010011111101: color_data = 12'b001110100111;
		16'b0010010011111110: color_data = 12'b001110100111;
		16'b0010010011111111: color_data = 12'b001110100111;
		16'b0010010100000000: color_data = 12'b001110100111;
		16'b0010010100000001: color_data = 12'b001110100111;
		16'b0010010100000010: color_data = 12'b001110100111;
		16'b0010010100000011: color_data = 12'b001110100111;
		16'b0010010100000100: color_data = 12'b001110100111;
		16'b0010010100000101: color_data = 12'b001110100111;
		16'b0010010100000110: color_data = 12'b001110100111;
		16'b0010010100000111: color_data = 12'b001110100111;
		16'b0010010100001000: color_data = 12'b001110100111;
		16'b0010010100001001: color_data = 12'b001110100111;
		16'b0010010100001010: color_data = 12'b001110100111;
		16'b0010010100001011: color_data = 12'b001110100111;
		16'b0010010100001100: color_data = 12'b001110100111;
		16'b0010010100001101: color_data = 12'b001110100111;
		16'b0010010100001110: color_data = 12'b001110100111;
		16'b0010010100001111: color_data = 12'b001110100111;
		16'b0010010100010000: color_data = 12'b001110100111;
		16'b0010010100010001: color_data = 12'b001110100111;
		16'b0010010100010010: color_data = 12'b001110100111;
		16'b0010010100010011: color_data = 12'b001110100111;
		16'b0010010100010100: color_data = 12'b001110100111;
		16'b0010010100010101: color_data = 12'b001110100111;
		16'b0010010100010110: color_data = 12'b001110100111;
		16'b0010010100010111: color_data = 12'b001110100111;
		16'b0010010100011000: color_data = 12'b001110100111;
		16'b0010010100011001: color_data = 12'b001110100111;
		16'b0010010100011010: color_data = 12'b001110100111;
		16'b0010010100011011: color_data = 12'b001110100111;
		16'b0010010100011100: color_data = 12'b001110100111;
		16'b0010010100011101: color_data = 12'b001110100111;
		16'b0010010100011110: color_data = 12'b001110100111;
		16'b0010010100011111: color_data = 12'b001110100111;
		16'b0010010100100000: color_data = 12'b001110100111;
		16'b0010010100100001: color_data = 12'b001110100111;
		16'b0010010100100010: color_data = 12'b001110100111;
		16'b0010010100100011: color_data = 12'b001110100111;
		16'b0010010100100100: color_data = 12'b001110100111;
		16'b0010010100100101: color_data = 12'b001110100111;
		16'b0010010100100110: color_data = 12'b001110100111;
		16'b0010010100101101: color_data = 12'b001110100111;
		16'b0010010100101110: color_data = 12'b001110100111;
		16'b0010010100101111: color_data = 12'b001110100111;
		16'b0010010100110000: color_data = 12'b001110100111;
		16'b0010010100110001: color_data = 12'b001110100111;
		16'b0010010100110010: color_data = 12'b001110100111;
		16'b0010010100110011: color_data = 12'b001110100111;
		16'b0010010100110100: color_data = 12'b001110100111;
		16'b0010010100110101: color_data = 12'b001110100111;
		16'b0010010100110110: color_data = 12'b001110100111;
		16'b0010010100110111: color_data = 12'b001110100111;
		16'b0010010100111000: color_data = 12'b001110100111;
		16'b0010010100111001: color_data = 12'b001110100111;
		16'b0010010100111010: color_data = 12'b001110100111;
		16'b0010010100111011: color_data = 12'b001110100111;
		16'b0010010100111100: color_data = 12'b001110100111;
		16'b0010010100111101: color_data = 12'b001110100111;
		16'b0010010100111110: color_data = 12'b001110100111;
		16'b0010010100111111: color_data = 12'b001110100111;
		16'b0010010101000000: color_data = 12'b001110100111;
		16'b0010010101000001: color_data = 12'b001110100111;
		16'b0010010101000010: color_data = 12'b001110100111;
		16'b0010010101000011: color_data = 12'b001110100111;
		16'b0010010101000100: color_data = 12'b001110100111;
		16'b0010010101000101: color_data = 12'b001110100111;
		16'b0010010101000110: color_data = 12'b001110100111;
		16'b0010010101000111: color_data = 12'b001110100111;
		16'b0010010101001000: color_data = 12'b001110100111;
		16'b0010010101001001: color_data = 12'b001110100111;
		16'b0010010101001010: color_data = 12'b001110100111;
		16'b0010010101011110: color_data = 12'b001110100111;
		16'b0010010101011111: color_data = 12'b001110100111;
		16'b0010010101100000: color_data = 12'b001110100111;
		16'b0010010101100001: color_data = 12'b001110100111;
		16'b0010010101100010: color_data = 12'b001110100111;
		16'b0010010101100011: color_data = 12'b001110100111;
		16'b0010010101100100: color_data = 12'b001110100111;
		16'b0010010101100101: color_data = 12'b001110100111;
		16'b0010010101100110: color_data = 12'b001110100111;
		16'b0010010101100111: color_data = 12'b001110100111;
		16'b0010010101101000: color_data = 12'b001110100111;
		16'b0010010101101001: color_data = 12'b001110100111;
		16'b0010010101101010: color_data = 12'b001110100111;
		16'b0010010101101011: color_data = 12'b001110100111;
		16'b0010010101101100: color_data = 12'b001110100111;
		16'b0010010101101101: color_data = 12'b001110100111;
		16'b0010010101101110: color_data = 12'b001110100111;
		16'b0010010101101111: color_data = 12'b001110100111;
		16'b0010010101110000: color_data = 12'b001110100111;
		16'b0010010101110001: color_data = 12'b001110100111;
		16'b0010010101110010: color_data = 12'b001110100111;
		16'b0010010101110011: color_data = 12'b001110100111;
		16'b0010010101110100: color_data = 12'b001110100111;
		16'b0010010101110101: color_data = 12'b001110100111;
		16'b0010010101110110: color_data = 12'b001110100111;
		16'b0010010101110111: color_data = 12'b001110100111;
		16'b0010010101111000: color_data = 12'b001110100111;
		16'b0010010101111001: color_data = 12'b001110100111;
		16'b0010010101111010: color_data = 12'b001110100111;
		16'b0010010101111011: color_data = 12'b001110100111;
		16'b0010011000000111: color_data = 12'b001110100111;
		16'b0010011000001000: color_data = 12'b001110100111;
		16'b0010011000001001: color_data = 12'b001110100111;
		16'b0010011000001010: color_data = 12'b001110100111;
		16'b0010011000001011: color_data = 12'b001110100111;
		16'b0010011000001100: color_data = 12'b001110100111;
		16'b0010011000001101: color_data = 12'b001110100111;
		16'b0010011000001110: color_data = 12'b001110100111;
		16'b0010011000001111: color_data = 12'b001110100111;
		16'b0010011000010000: color_data = 12'b001110100111;
		16'b0010011000010001: color_data = 12'b001110100111;
		16'b0010011000010010: color_data = 12'b001110100111;
		16'b0010011000010011: color_data = 12'b001110100111;
		16'b0010011000010100: color_data = 12'b001110100111;
		16'b0010011000010101: color_data = 12'b001110100111;
		16'b0010011000010110: color_data = 12'b001110100111;
		16'b0010011000010111: color_data = 12'b001110100111;
		16'b0010011000011000: color_data = 12'b001110100111;
		16'b0010011000011001: color_data = 12'b001110100111;
		16'b0010011000011010: color_data = 12'b001110100111;
		16'b0010011000011011: color_data = 12'b001110100111;
		16'b0010011000011100: color_data = 12'b001110100111;
		16'b0010011000011101: color_data = 12'b001110100111;
		16'b0010011000011110: color_data = 12'b001110100111;
		16'b0010011000011111: color_data = 12'b001110100111;
		16'b0010011000100000: color_data = 12'b001110100111;
		16'b0010011000100001: color_data = 12'b001110100111;
		16'b0010011000100010: color_data = 12'b001110100111;
		16'b0010011000100011: color_data = 12'b001110100111;
		16'b0010011000100100: color_data = 12'b001110100111;
		16'b0010011000101011: color_data = 12'b001110100111;
		16'b0010011000101100: color_data = 12'b001110100111;
		16'b0010011000101101: color_data = 12'b001110100111;
		16'b0010011000101110: color_data = 12'b001110100111;
		16'b0010011000101111: color_data = 12'b001110100111;
		16'b0010011000110000: color_data = 12'b001110100111;
		16'b0010011000110001: color_data = 12'b001110100111;
		16'b0010011000110010: color_data = 12'b001110100111;
		16'b0010011000110011: color_data = 12'b001110100111;
		16'b0010011000110100: color_data = 12'b001110100111;
		16'b0010011000110101: color_data = 12'b001110100111;
		16'b0010011000110110: color_data = 12'b001110100111;
		16'b0010011000110111: color_data = 12'b001110100111;
		16'b0010011001000100: color_data = 12'b001110100111;
		16'b0010011001000101: color_data = 12'b001110100111;
		16'b0010011001000110: color_data = 12'b001110100111;
		16'b0010011001000111: color_data = 12'b001110100111;
		16'b0010011001001000: color_data = 12'b001110100111;
		16'b0010011001001001: color_data = 12'b001110100111;
		16'b0010011001001010: color_data = 12'b001110100111;
		16'b0010011001001011: color_data = 12'b001110100111;
		16'b0010011001001100: color_data = 12'b001110100111;
		16'b0010011001001101: color_data = 12'b001110100111;
		16'b0010011001001110: color_data = 12'b001110100111;
		16'b0010011001001111: color_data = 12'b001110100111;
		16'b0010011001010110: color_data = 12'b001110100111;
		16'b0010011001010111: color_data = 12'b001110100111;
		16'b0010011001011000: color_data = 12'b001110100111;
		16'b0010011001011001: color_data = 12'b001110100111;
		16'b0010011001011010: color_data = 12'b001110100111;
		16'b0010011001011011: color_data = 12'b001110100111;
		16'b0010011001011100: color_data = 12'b001110100111;
		16'b0010011001011101: color_data = 12'b001110100111;
		16'b0010011001011110: color_data = 12'b001110100111;
		16'b0010011001011111: color_data = 12'b001110100111;
		16'b0010011001100000: color_data = 12'b001110100111;
		16'b0010011001100001: color_data = 12'b001110100111;
		16'b0010011001100010: color_data = 12'b001110100111;
		16'b0010011001100011: color_data = 12'b001110100111;
		16'b0010011001100100: color_data = 12'b001110100111;
		16'b0010011001100101: color_data = 12'b001110100111;
		16'b0010011001100110: color_data = 12'b001110100111;
		16'b0010011001100111: color_data = 12'b001110100111;
		16'b0010011001101000: color_data = 12'b001110100111;
		16'b0010011001101001: color_data = 12'b001110100111;
		16'b0010011001101010: color_data = 12'b001110100111;
		16'b0010011001101011: color_data = 12'b001110100111;
		16'b0010011001101100: color_data = 12'b001110100111;
		16'b0010011001101101: color_data = 12'b001110100111;
		16'b0010011001101110: color_data = 12'b001110100111;
		16'b0010011001110101: color_data = 12'b001110100111;
		16'b0010011001110110: color_data = 12'b001110100111;
		16'b0010011001110111: color_data = 12'b001110100111;
		16'b0010011001111000: color_data = 12'b001110100111;
		16'b0010011001111001: color_data = 12'b001110100111;
		16'b0010011001111010: color_data = 12'b001110100111;
		16'b0010011001111011: color_data = 12'b001110100111;
		16'b0010011001111100: color_data = 12'b001110100111;
		16'b0010011001111101: color_data = 12'b001110100111;
		16'b0010011001111110: color_data = 12'b001110100111;
		16'b0010011001111111: color_data = 12'b001110100111;
		16'b0010011010000000: color_data = 12'b001110100111;
		16'b0010011010000001: color_data = 12'b001110100111;
		16'b0010011010000010: color_data = 12'b001110100111;
		16'b0010011010000011: color_data = 12'b001110100111;
		16'b0010011010000100: color_data = 12'b001110100111;
		16'b0010011010000101: color_data = 12'b001110100111;
		16'b0010011010000110: color_data = 12'b001110100111;
		16'b0010011010000111: color_data = 12'b001110100111;
		16'b0010011010001000: color_data = 12'b001110100111;
		16'b0010011010001001: color_data = 12'b001110100111;
		16'b0010011010001010: color_data = 12'b001110100111;
		16'b0010011010001011: color_data = 12'b001110100111;
		16'b0010011010001100: color_data = 12'b001110100111;
		16'b0010011010001101: color_data = 12'b001110100111;
		16'b0010011010001110: color_data = 12'b001110100111;
		16'b0010011010001111: color_data = 12'b001110100111;
		16'b0010011010010000: color_data = 12'b001110100111;
		16'b0010011010010001: color_data = 12'b001110100111;
		16'b0010011010010010: color_data = 12'b001110100111;
		16'b0010011010010011: color_data = 12'b001110100111;
		16'b0010011010100110: color_data = 12'b001110100111;
		16'b0010011010100111: color_data = 12'b001110100111;
		16'b0010011010101000: color_data = 12'b001110100111;
		16'b0010011010101001: color_data = 12'b001110100111;
		16'b0010011010101010: color_data = 12'b001110100111;
		16'b0010011010101011: color_data = 12'b001110100111;
		16'b0010011010101100: color_data = 12'b001110100111;
		16'b0010011010101101: color_data = 12'b001110100111;
		16'b0010011010101110: color_data = 12'b001110100111;
		16'b0010011010101111: color_data = 12'b001110100111;
		16'b0010011010110000: color_data = 12'b001110100111;
		16'b0010011010110001: color_data = 12'b001110100111;
		16'b0010011010110010: color_data = 12'b001110100111;
		16'b0010011010110011: color_data = 12'b001110100111;
		16'b0010011010110100: color_data = 12'b001110100111;
		16'b0010011010110101: color_data = 12'b001110100111;
		16'b0010011010110110: color_data = 12'b001110100111;
		16'b0010011010110111: color_data = 12'b001110100111;
		16'b0010011010111000: color_data = 12'b001110100111;
		16'b0010011010111001: color_data = 12'b001110100111;
		16'b0010011010111010: color_data = 12'b001110100111;
		16'b0010011010111011: color_data = 12'b001110100111;
		16'b0010011010111100: color_data = 12'b001110100111;
		16'b0010011010111101: color_data = 12'b001110100111;
		16'b0010011010111110: color_data = 12'b001110100111;
		16'b0010011010111111: color_data = 12'b001110100111;
		16'b0010011011000000: color_data = 12'b001110100111;
		16'b0010011011000001: color_data = 12'b001110100111;
		16'b0010011011000010: color_data = 12'b001110100111;
		16'b0010011011000011: color_data = 12'b001110100111;
		16'b0010011011000100: color_data = 12'b001110100111;
		16'b0010011011001011: color_data = 12'b001110100111;
		16'b0010011011001100: color_data = 12'b001110100111;
		16'b0010011011001101: color_data = 12'b001110100111;
		16'b0010011011001110: color_data = 12'b001110100111;
		16'b0010011011001111: color_data = 12'b001110100111;
		16'b0010011011010000: color_data = 12'b001110100111;
		16'b0010011011010001: color_data = 12'b001110100111;
		16'b0010011011010010: color_data = 12'b001110100111;
		16'b0010011011010011: color_data = 12'b001110100111;
		16'b0010011011010100: color_data = 12'b001110100111;
		16'b0010011011010101: color_data = 12'b001110100111;
		16'b0010011011010110: color_data = 12'b001110100111;
		16'b0010011011010111: color_data = 12'b001110100111;
		16'b0010011011011000: color_data = 12'b001110100111;
		16'b0010011011011001: color_data = 12'b001110100111;
		16'b0010011011011010: color_data = 12'b001110100111;
		16'b0010011011011011: color_data = 12'b001110100111;
		16'b0010011011011100: color_data = 12'b001110100111;
		16'b0010011011011101: color_data = 12'b001110100111;
		16'b0010011011011110: color_data = 12'b001110100111;
		16'b0010011011011111: color_data = 12'b001110100111;
		16'b0010011011100000: color_data = 12'b001110100111;
		16'b0010011011100001: color_data = 12'b001110100111;
		16'b0010011011100010: color_data = 12'b001110100111;
		16'b0010011011100011: color_data = 12'b001110100111;
		16'b0010011011100100: color_data = 12'b001110100111;
		16'b0010011011100101: color_data = 12'b001110100111;
		16'b0010011011100110: color_data = 12'b001110100111;
		16'b0010011011100111: color_data = 12'b001110100111;
		16'b0010011011101000: color_data = 12'b001110100111;
		16'b0010011011101001: color_data = 12'b001110100111;
		16'b0010011011101010: color_data = 12'b001110100111;
		16'b0010011011101011: color_data = 12'b001110100111;
		16'b0010011011101100: color_data = 12'b001110100111;
		16'b0010011011101101: color_data = 12'b001110100111;
		16'b0010011011101110: color_data = 12'b001110100111;
		16'b0010011011101111: color_data = 12'b001110100111;
		16'b0010011011110110: color_data = 12'b001110100111;
		16'b0010011011110111: color_data = 12'b001110100111;
		16'b0010011011111000: color_data = 12'b001110100111;
		16'b0010011011111001: color_data = 12'b001110100111;
		16'b0010011011111010: color_data = 12'b001110100111;
		16'b0010011011111011: color_data = 12'b001110100111;
		16'b0010011011111100: color_data = 12'b001110100111;
		16'b0010011011111101: color_data = 12'b001110100111;
		16'b0010011011111110: color_data = 12'b001110100111;
		16'b0010011011111111: color_data = 12'b001110100111;
		16'b0010011100000000: color_data = 12'b001110100111;
		16'b0010011100000001: color_data = 12'b001110100111;
		16'b0010011100000010: color_data = 12'b001110100111;
		16'b0010011100000011: color_data = 12'b001110100111;
		16'b0010011100000100: color_data = 12'b001110100111;
		16'b0010011100000101: color_data = 12'b001110100111;
		16'b0010011100000110: color_data = 12'b001110100111;
		16'b0010011100000111: color_data = 12'b001110100111;
		16'b0010011100001000: color_data = 12'b001110100111;
		16'b0010011100001001: color_data = 12'b001110100111;
		16'b0010011100001010: color_data = 12'b001110100111;
		16'b0010011100001011: color_data = 12'b001110100111;
		16'b0010011100001100: color_data = 12'b001110100111;
		16'b0010011100001101: color_data = 12'b001110100111;
		16'b0010011100001110: color_data = 12'b001110100111;
		16'b0010011100001111: color_data = 12'b001110100111;
		16'b0010011100010000: color_data = 12'b001110100111;
		16'b0010011100010001: color_data = 12'b001110100111;
		16'b0010011100010010: color_data = 12'b001110100111;
		16'b0010011100010011: color_data = 12'b001110100111;
		16'b0010011100010100: color_data = 12'b001110100111;
		16'b0010011100010101: color_data = 12'b001110100111;
		16'b0010011100010110: color_data = 12'b001110100111;
		16'b0010011100010111: color_data = 12'b001110100111;
		16'b0010011100011000: color_data = 12'b001110100111;
		16'b0010011100011001: color_data = 12'b001110100111;
		16'b0010011100011010: color_data = 12'b001110100111;
		16'b0010011100011011: color_data = 12'b001110100111;
		16'b0010011100011100: color_data = 12'b001110100111;
		16'b0010011100011101: color_data = 12'b001110100111;
		16'b0010011100011110: color_data = 12'b001110100111;
		16'b0010011100011111: color_data = 12'b001110100111;
		16'b0010011100100000: color_data = 12'b001110100111;
		16'b0010011100100001: color_data = 12'b001110100111;
		16'b0010011100100010: color_data = 12'b001110100111;
		16'b0010011100100011: color_data = 12'b001110100111;
		16'b0010011100100100: color_data = 12'b001110100111;
		16'b0010011100100101: color_data = 12'b001110100111;
		16'b0010011100100110: color_data = 12'b001110100111;
		16'b0010011100101101: color_data = 12'b001110100111;
		16'b0010011100101110: color_data = 12'b001110100111;
		16'b0010011100101111: color_data = 12'b001110100111;
		16'b0010011100110000: color_data = 12'b001110100111;
		16'b0010011100110001: color_data = 12'b001110100111;
		16'b0010011100110010: color_data = 12'b001110100111;
		16'b0010011100110011: color_data = 12'b001110100111;
		16'b0010011100110100: color_data = 12'b001110100111;
		16'b0010011100110101: color_data = 12'b001110100111;
		16'b0010011100110110: color_data = 12'b001110100111;
		16'b0010011100110111: color_data = 12'b001110100111;
		16'b0010011100111000: color_data = 12'b001110100111;
		16'b0010011100111001: color_data = 12'b001110100111;
		16'b0010011100111010: color_data = 12'b001110100111;
		16'b0010011100111011: color_data = 12'b001110100111;
		16'b0010011100111100: color_data = 12'b001110100111;
		16'b0010011100111101: color_data = 12'b001110100111;
		16'b0010011100111110: color_data = 12'b001110100111;
		16'b0010011100111111: color_data = 12'b001110100111;
		16'b0010011101000000: color_data = 12'b001110100111;
		16'b0010011101000001: color_data = 12'b001110100111;
		16'b0010011101000010: color_data = 12'b001110100111;
		16'b0010011101000011: color_data = 12'b001110100111;
		16'b0010011101000100: color_data = 12'b001110100111;
		16'b0010011101000101: color_data = 12'b001110100111;
		16'b0010011101000110: color_data = 12'b001110100111;
		16'b0010011101000111: color_data = 12'b001110100111;
		16'b0010011101001000: color_data = 12'b001110100111;
		16'b0010011101001001: color_data = 12'b001110100111;
		16'b0010011101001010: color_data = 12'b001110100111;
		16'b0010011101011110: color_data = 12'b001110100111;
		16'b0010011101011111: color_data = 12'b001110100111;
		16'b0010011101100000: color_data = 12'b001110100111;
		16'b0010011101100001: color_data = 12'b001110100111;
		16'b0010011101100010: color_data = 12'b001110100111;
		16'b0010011101100011: color_data = 12'b001110100111;
		16'b0010011101100100: color_data = 12'b001110100111;
		16'b0010011101100101: color_data = 12'b001110100111;
		16'b0010011101100110: color_data = 12'b001110100111;
		16'b0010011101100111: color_data = 12'b001110100111;
		16'b0010011101101000: color_data = 12'b001110100111;
		16'b0010011101101001: color_data = 12'b001110100111;
		16'b0010011101101010: color_data = 12'b001110100111;
		16'b0010011101101011: color_data = 12'b001110100111;
		16'b0010011101101100: color_data = 12'b001110100111;
		16'b0010011101101101: color_data = 12'b001110100111;
		16'b0010011101101110: color_data = 12'b001110100111;
		16'b0010011101101111: color_data = 12'b001110100111;
		16'b0010011101110000: color_data = 12'b001110100111;
		16'b0010011101110001: color_data = 12'b001110100111;
		16'b0010011101110010: color_data = 12'b001110100111;
		16'b0010011101110011: color_data = 12'b001110100111;
		16'b0010011101110100: color_data = 12'b001110100111;
		16'b0010011101110101: color_data = 12'b001110100111;
		16'b0010011101110110: color_data = 12'b001110100111;
		16'b0010011101110111: color_data = 12'b001110100111;
		16'b0010011101111000: color_data = 12'b001110100111;
		16'b0010011101111001: color_data = 12'b001110100111;
		16'b0010011101111010: color_data = 12'b001110100111;
		16'b0010011101111011: color_data = 12'b001110100111;
		16'b0010100000000111: color_data = 12'b001110100111;
		16'b0010100000001000: color_data = 12'b001110100111;
		16'b0010100000001001: color_data = 12'b001110100111;
		16'b0010100000001010: color_data = 12'b001110100111;
		16'b0010100000001011: color_data = 12'b001110100111;
		16'b0010100000001100: color_data = 12'b001110100111;
		16'b0010100000001101: color_data = 12'b001110100111;
		16'b0010100000001110: color_data = 12'b001110100111;
		16'b0010100000001111: color_data = 12'b001110100111;
		16'b0010100000010000: color_data = 12'b001110100111;
		16'b0010100000010001: color_data = 12'b001110100111;
		16'b0010100000010010: color_data = 12'b001110100111;
		16'b0010100000010011: color_data = 12'b001110100111;
		16'b0010100000010100: color_data = 12'b001110100111;
		16'b0010100000010101: color_data = 12'b001110100111;
		16'b0010100000010110: color_data = 12'b001110100111;
		16'b0010100000010111: color_data = 12'b001110100111;
		16'b0010100000011000: color_data = 12'b001110100111;
		16'b0010100000011001: color_data = 12'b001110100111;
		16'b0010100000011010: color_data = 12'b001110100111;
		16'b0010100000011011: color_data = 12'b001110100111;
		16'b0010100000011100: color_data = 12'b001110100111;
		16'b0010100000011101: color_data = 12'b001110100111;
		16'b0010100000011110: color_data = 12'b001110100111;
		16'b0010100000011111: color_data = 12'b001110100111;
		16'b0010100000100000: color_data = 12'b001110100111;
		16'b0010100000100001: color_data = 12'b001110100111;
		16'b0010100000100010: color_data = 12'b001110100111;
		16'b0010100000100011: color_data = 12'b001110100111;
		16'b0010100000100100: color_data = 12'b001110100111;
		16'b0010100000101011: color_data = 12'b001110100111;
		16'b0010100000101100: color_data = 12'b001110100111;
		16'b0010100000101101: color_data = 12'b001110100111;
		16'b0010100000101110: color_data = 12'b001110100111;
		16'b0010100000101111: color_data = 12'b001110100111;
		16'b0010100000110000: color_data = 12'b001110100111;
		16'b0010100000110001: color_data = 12'b001110100111;
		16'b0010100000110010: color_data = 12'b001110100111;
		16'b0010100000110011: color_data = 12'b001110100111;
		16'b0010100000110100: color_data = 12'b001110100111;
		16'b0010100000110101: color_data = 12'b001110100111;
		16'b0010100000110110: color_data = 12'b001110100111;
		16'b0010100000110111: color_data = 12'b001110100111;
		16'b0010100001000100: color_data = 12'b001110100111;
		16'b0010100001000101: color_data = 12'b001110100111;
		16'b0010100001000110: color_data = 12'b001110100111;
		16'b0010100001000111: color_data = 12'b001110100111;
		16'b0010100001001000: color_data = 12'b001110100111;
		16'b0010100001001001: color_data = 12'b001110100111;
		16'b0010100001001010: color_data = 12'b001110100111;
		16'b0010100001001011: color_data = 12'b001110100111;
		16'b0010100001001100: color_data = 12'b001110100111;
		16'b0010100001001101: color_data = 12'b001110100111;
		16'b0010100001001110: color_data = 12'b001110100111;
		16'b0010100001001111: color_data = 12'b001110100111;
		16'b0010100001010110: color_data = 12'b001110100111;
		16'b0010100001010111: color_data = 12'b001110100111;
		16'b0010100001011000: color_data = 12'b001110100111;
		16'b0010100001011001: color_data = 12'b001110100111;
		16'b0010100001011010: color_data = 12'b001110100111;
		16'b0010100001011011: color_data = 12'b001110100111;
		16'b0010100001011100: color_data = 12'b001110100111;
		16'b0010100001011101: color_data = 12'b001110100111;
		16'b0010100001011110: color_data = 12'b001110100111;
		16'b0010100001011111: color_data = 12'b001110100111;
		16'b0010100001100000: color_data = 12'b001110100111;
		16'b0010100001100001: color_data = 12'b001110100111;
		16'b0010100001100010: color_data = 12'b001110100111;
		16'b0010100001100011: color_data = 12'b001110100111;
		16'b0010100001100100: color_data = 12'b001110100111;
		16'b0010100001100101: color_data = 12'b001110100111;
		16'b0010100001100110: color_data = 12'b001110100111;
		16'b0010100001100111: color_data = 12'b001110100111;
		16'b0010100001101000: color_data = 12'b001110100111;
		16'b0010100001101001: color_data = 12'b001110100111;
		16'b0010100001101010: color_data = 12'b001110100111;
		16'b0010100001101011: color_data = 12'b001110100111;
		16'b0010100001101100: color_data = 12'b001110100111;
		16'b0010100001101101: color_data = 12'b001110100111;
		16'b0010100001101110: color_data = 12'b001110100111;
		16'b0010100001110101: color_data = 12'b001110100111;
		16'b0010100001110110: color_data = 12'b001110100111;
		16'b0010100001110111: color_data = 12'b001110100111;
		16'b0010100001111000: color_data = 12'b001110100111;
		16'b0010100001111001: color_data = 12'b001110100111;
		16'b0010100001111010: color_data = 12'b001110100111;
		16'b0010100001111011: color_data = 12'b001110100111;
		16'b0010100001111100: color_data = 12'b001110100111;
		16'b0010100001111101: color_data = 12'b001110100111;
		16'b0010100001111110: color_data = 12'b001110100111;
		16'b0010100001111111: color_data = 12'b001110100111;
		16'b0010100010000000: color_data = 12'b001110100111;
		16'b0010100010000001: color_data = 12'b001110100111;
		16'b0010100010000010: color_data = 12'b001110100111;
		16'b0010100010000011: color_data = 12'b001110100111;
		16'b0010100010000100: color_data = 12'b001110100111;
		16'b0010100010000101: color_data = 12'b001110100111;
		16'b0010100010000110: color_data = 12'b001110100111;
		16'b0010100010000111: color_data = 12'b001110100111;
		16'b0010100010001000: color_data = 12'b001110100111;
		16'b0010100010001001: color_data = 12'b001110100111;
		16'b0010100010001010: color_data = 12'b001110100111;
		16'b0010100010001011: color_data = 12'b001110100111;
		16'b0010100010001100: color_data = 12'b001110100111;
		16'b0010100010001101: color_data = 12'b001110100111;
		16'b0010100010001110: color_data = 12'b001110100111;
		16'b0010100010001111: color_data = 12'b001110100111;
		16'b0010100010010000: color_data = 12'b001110100111;
		16'b0010100010010001: color_data = 12'b001110100111;
		16'b0010100010010010: color_data = 12'b001110100111;
		16'b0010100010010011: color_data = 12'b001110100111;
		16'b0010100010100110: color_data = 12'b001110100111;
		16'b0010100010100111: color_data = 12'b001110100111;
		16'b0010100010101000: color_data = 12'b001110100111;
		16'b0010100010101001: color_data = 12'b001110100111;
		16'b0010100010101010: color_data = 12'b001110100111;
		16'b0010100010101011: color_data = 12'b001110100111;
		16'b0010100010101100: color_data = 12'b001110100111;
		16'b0010100010101101: color_data = 12'b001110100111;
		16'b0010100010101110: color_data = 12'b001110100111;
		16'b0010100010101111: color_data = 12'b001110100111;
		16'b0010100010110000: color_data = 12'b001110100111;
		16'b0010100010110001: color_data = 12'b001110100111;
		16'b0010100010110010: color_data = 12'b001110100111;
		16'b0010100010110011: color_data = 12'b001110100111;
		16'b0010100010110100: color_data = 12'b001110100111;
		16'b0010100010110101: color_data = 12'b001110100111;
		16'b0010100010110110: color_data = 12'b001110100111;
		16'b0010100010110111: color_data = 12'b001110100111;
		16'b0010100010111000: color_data = 12'b001110100111;
		16'b0010100010111001: color_data = 12'b001110100111;
		16'b0010100010111010: color_data = 12'b001110100111;
		16'b0010100010111011: color_data = 12'b001110100111;
		16'b0010100010111100: color_data = 12'b001110100111;
		16'b0010100010111101: color_data = 12'b001110100111;
		16'b0010100010111110: color_data = 12'b001110100111;
		16'b0010100010111111: color_data = 12'b001110100111;
		16'b0010100011000000: color_data = 12'b001110100111;
		16'b0010100011000001: color_data = 12'b001110100111;
		16'b0010100011000010: color_data = 12'b001110100111;
		16'b0010100011000011: color_data = 12'b001110100111;
		16'b0010100011000100: color_data = 12'b001110100111;
		16'b0010100011001011: color_data = 12'b001110100111;
		16'b0010100011001100: color_data = 12'b001110100111;
		16'b0010100011001101: color_data = 12'b001110100111;
		16'b0010100011001110: color_data = 12'b001110100111;
		16'b0010100011001111: color_data = 12'b001110100111;
		16'b0010100011010000: color_data = 12'b001110100111;
		16'b0010100011010001: color_data = 12'b001110100111;
		16'b0010100011010010: color_data = 12'b001110100111;
		16'b0010100011010011: color_data = 12'b001110100111;
		16'b0010100011010100: color_data = 12'b001110100111;
		16'b0010100011010101: color_data = 12'b001110100111;
		16'b0010100011010110: color_data = 12'b001110100111;
		16'b0010100011010111: color_data = 12'b001110100111;
		16'b0010100011011000: color_data = 12'b001110100111;
		16'b0010100011011001: color_data = 12'b001110100111;
		16'b0010100011011010: color_data = 12'b001110100111;
		16'b0010100011011011: color_data = 12'b001110100111;
		16'b0010100011011100: color_data = 12'b001110100111;
		16'b0010100011011101: color_data = 12'b001110100111;
		16'b0010100011011110: color_data = 12'b001110100111;
		16'b0010100011011111: color_data = 12'b001110100111;
		16'b0010100011100000: color_data = 12'b001110100111;
		16'b0010100011100001: color_data = 12'b001110100111;
		16'b0010100011100010: color_data = 12'b001110100111;
		16'b0010100011100011: color_data = 12'b001110100111;
		16'b0010100011100100: color_data = 12'b001110100111;
		16'b0010100011100101: color_data = 12'b001110100111;
		16'b0010100011100110: color_data = 12'b001110100111;
		16'b0010100011100111: color_data = 12'b001110100111;
		16'b0010100011101000: color_data = 12'b001110100111;
		16'b0010100011101001: color_data = 12'b001110100111;
		16'b0010100011101010: color_data = 12'b001110100111;
		16'b0010100011101011: color_data = 12'b001110100111;
		16'b0010100011101100: color_data = 12'b001110100111;
		16'b0010100011101101: color_data = 12'b001110100111;
		16'b0010100011101110: color_data = 12'b001110100111;
		16'b0010100011101111: color_data = 12'b001110100111;
		16'b0010100011110110: color_data = 12'b001110100111;
		16'b0010100011110111: color_data = 12'b001110100111;
		16'b0010100011111000: color_data = 12'b001110100111;
		16'b0010100011111001: color_data = 12'b001110100111;
		16'b0010100011111010: color_data = 12'b001110100111;
		16'b0010100011111011: color_data = 12'b001110100111;
		16'b0010100011111100: color_data = 12'b001110100111;
		16'b0010100011111101: color_data = 12'b001110100111;
		16'b0010100011111110: color_data = 12'b001110100111;
		16'b0010100011111111: color_data = 12'b001110100111;
		16'b0010100100000000: color_data = 12'b001110100111;
		16'b0010100100000001: color_data = 12'b001110100111;
		16'b0010100100000010: color_data = 12'b001110100111;
		16'b0010100100000011: color_data = 12'b001110100111;
		16'b0010100100000100: color_data = 12'b001110100111;
		16'b0010100100000101: color_data = 12'b001110100111;
		16'b0010100100000110: color_data = 12'b001110100111;
		16'b0010100100000111: color_data = 12'b001110100111;
		16'b0010100100001000: color_data = 12'b001110100111;
		16'b0010100100001001: color_data = 12'b001110100111;
		16'b0010100100001010: color_data = 12'b001110100111;
		16'b0010100100001011: color_data = 12'b001110100111;
		16'b0010100100001100: color_data = 12'b001110100111;
		16'b0010100100001101: color_data = 12'b001110100111;
		16'b0010100100001110: color_data = 12'b001110100111;
		16'b0010100100001111: color_data = 12'b001110100111;
		16'b0010100100010000: color_data = 12'b001110100111;
		16'b0010100100010001: color_data = 12'b001110100111;
		16'b0010100100010010: color_data = 12'b001110100111;
		16'b0010100100010011: color_data = 12'b001110100111;
		16'b0010100100010100: color_data = 12'b001110100111;
		16'b0010100100010101: color_data = 12'b001110100111;
		16'b0010100100010110: color_data = 12'b001110100111;
		16'b0010100100010111: color_data = 12'b001110100111;
		16'b0010100100011000: color_data = 12'b001110100111;
		16'b0010100100011001: color_data = 12'b001110100111;
		16'b0010100100011010: color_data = 12'b001110100111;
		16'b0010100100011011: color_data = 12'b001110100111;
		16'b0010100100011100: color_data = 12'b001110100111;
		16'b0010100100011101: color_data = 12'b001110100111;
		16'b0010100100011110: color_data = 12'b001110100111;
		16'b0010100100011111: color_data = 12'b001110100111;
		16'b0010100100100000: color_data = 12'b001110100111;
		16'b0010100100100001: color_data = 12'b001110100111;
		16'b0010100100100010: color_data = 12'b001110100111;
		16'b0010100100100011: color_data = 12'b001110100111;
		16'b0010100100100100: color_data = 12'b001110100111;
		16'b0010100100100101: color_data = 12'b001110100111;
		16'b0010100100100110: color_data = 12'b001110100111;
		16'b0010100100101101: color_data = 12'b001110100111;
		16'b0010100100101110: color_data = 12'b001110100111;
		16'b0010100100101111: color_data = 12'b001110100111;
		16'b0010100100110000: color_data = 12'b001110100111;
		16'b0010100100110001: color_data = 12'b001110100111;
		16'b0010100100110010: color_data = 12'b001110100111;
		16'b0010100100110011: color_data = 12'b001110100111;
		16'b0010100100110100: color_data = 12'b001110100111;
		16'b0010100100110101: color_data = 12'b001110100111;
		16'b0010100100110110: color_data = 12'b001110100111;
		16'b0010100100110111: color_data = 12'b001110100111;
		16'b0010100100111000: color_data = 12'b001110100111;
		16'b0010100100111001: color_data = 12'b001110100111;
		16'b0010100100111010: color_data = 12'b001110100111;
		16'b0010100100111011: color_data = 12'b001110100111;
		16'b0010100100111100: color_data = 12'b001110100111;
		16'b0010100100111101: color_data = 12'b001110100111;
		16'b0010100100111110: color_data = 12'b001110100111;
		16'b0010100100111111: color_data = 12'b001110100111;
		16'b0010100101000000: color_data = 12'b001110100111;
		16'b0010100101000001: color_data = 12'b001110100111;
		16'b0010100101000010: color_data = 12'b001110100111;
		16'b0010100101000011: color_data = 12'b001110100111;
		16'b0010100101000100: color_data = 12'b001110100111;
		16'b0010100101000101: color_data = 12'b001110100111;
		16'b0010100101000110: color_data = 12'b001110100111;
		16'b0010100101000111: color_data = 12'b001110100111;
		16'b0010100101001000: color_data = 12'b001110100111;
		16'b0010100101001001: color_data = 12'b001110100111;
		16'b0010100101001010: color_data = 12'b001110100111;
		16'b0010100101011110: color_data = 12'b001110100111;
		16'b0010100101011111: color_data = 12'b001110100111;
		16'b0010100101100000: color_data = 12'b001110100111;
		16'b0010100101100001: color_data = 12'b001110100111;
		16'b0010100101100010: color_data = 12'b001110100111;
		16'b0010100101100011: color_data = 12'b001110100111;
		16'b0010100101100100: color_data = 12'b001110100111;
		16'b0010100101100101: color_data = 12'b001110100111;
		16'b0010100101100110: color_data = 12'b001110100111;
		16'b0010100101100111: color_data = 12'b001110100111;
		16'b0010100101101000: color_data = 12'b001110100111;
		16'b0010100101101001: color_data = 12'b001110100111;
		16'b0010100101101010: color_data = 12'b001110100111;
		16'b0010100101101011: color_data = 12'b001110100111;
		16'b0010100101101100: color_data = 12'b001110100111;
		16'b0010100101101101: color_data = 12'b001110100111;
		16'b0010100101101110: color_data = 12'b001110100111;
		16'b0010100101101111: color_data = 12'b001110100111;
		16'b0010100101110000: color_data = 12'b001110100111;
		16'b0010100101110001: color_data = 12'b001110100111;
		16'b0010100101110010: color_data = 12'b001110100111;
		16'b0010100101110011: color_data = 12'b001110100111;
		16'b0010100101110100: color_data = 12'b001110100111;
		16'b0010100101110101: color_data = 12'b001110100111;
		16'b0010100101110110: color_data = 12'b001110100111;
		16'b0010100101110111: color_data = 12'b001110100111;
		16'b0010100101111000: color_data = 12'b001110100111;
		16'b0010100101111001: color_data = 12'b001110100111;
		16'b0010100101111010: color_data = 12'b001110100111;
		16'b0010100101111011: color_data = 12'b001110100111;
		16'b0010101000000111: color_data = 12'b001110100111;
		16'b0010101000001000: color_data = 12'b001110100111;
		16'b0010101000001001: color_data = 12'b001110100111;
		16'b0010101000001010: color_data = 12'b001110100111;
		16'b0010101000001011: color_data = 12'b001110100111;
		16'b0010101000001100: color_data = 12'b001110100111;
		16'b0010101000001101: color_data = 12'b001110100111;
		16'b0010101000001110: color_data = 12'b001110100111;
		16'b0010101000001111: color_data = 12'b001110100111;
		16'b0010101000010000: color_data = 12'b001110100111;
		16'b0010101000010001: color_data = 12'b001110100111;
		16'b0010101000010010: color_data = 12'b001110100111;
		16'b0010101000010011: color_data = 12'b001110100111;
		16'b0010101000010100: color_data = 12'b001110100111;
		16'b0010101000010101: color_data = 12'b001110100111;
		16'b0010101000010110: color_data = 12'b001110100111;
		16'b0010101000010111: color_data = 12'b001110100111;
		16'b0010101000011000: color_data = 12'b001110100111;
		16'b0010101000011001: color_data = 12'b001110100111;
		16'b0010101000011010: color_data = 12'b001110100111;
		16'b0010101000011011: color_data = 12'b001110100111;
		16'b0010101000011100: color_data = 12'b001110100111;
		16'b0010101000011101: color_data = 12'b001110100111;
		16'b0010101000011110: color_data = 12'b001110100111;
		16'b0010101000011111: color_data = 12'b001110100111;
		16'b0010101000100000: color_data = 12'b001110100111;
		16'b0010101000100001: color_data = 12'b001110100111;
		16'b0010101000100010: color_data = 12'b001110100111;
		16'b0010101000100011: color_data = 12'b001110100111;
		16'b0010101000100100: color_data = 12'b001110100111;
		16'b0010101000101011: color_data = 12'b001110100111;
		16'b0010101000101100: color_data = 12'b001110100111;
		16'b0010101000101101: color_data = 12'b001110100111;
		16'b0010101000101110: color_data = 12'b001110100111;
		16'b0010101000101111: color_data = 12'b001110100111;
		16'b0010101000110000: color_data = 12'b001110100111;
		16'b0010101000110001: color_data = 12'b001110100111;
		16'b0010101000110010: color_data = 12'b001110100111;
		16'b0010101000110011: color_data = 12'b001110100111;
		16'b0010101000110100: color_data = 12'b001110100111;
		16'b0010101000110101: color_data = 12'b001110100111;
		16'b0010101000110110: color_data = 12'b001110100111;
		16'b0010101000110111: color_data = 12'b001110100111;
		16'b0010101001000100: color_data = 12'b001110100111;
		16'b0010101001000101: color_data = 12'b001110100111;
		16'b0010101001000110: color_data = 12'b001110100111;
		16'b0010101001000111: color_data = 12'b001110100111;
		16'b0010101001001000: color_data = 12'b001110100111;
		16'b0010101001001001: color_data = 12'b001110100111;
		16'b0010101001001010: color_data = 12'b001110100111;
		16'b0010101001001011: color_data = 12'b001110100111;
		16'b0010101001001100: color_data = 12'b001110100111;
		16'b0010101001001101: color_data = 12'b001110100111;
		16'b0010101001001110: color_data = 12'b001110100111;
		16'b0010101001001111: color_data = 12'b001110100111;
		16'b0010101001010110: color_data = 12'b001110100111;
		16'b0010101001010111: color_data = 12'b001110100111;
		16'b0010101001011000: color_data = 12'b001110100111;
		16'b0010101001011001: color_data = 12'b001110100111;
		16'b0010101001011010: color_data = 12'b001110100111;
		16'b0010101001011011: color_data = 12'b001110100111;
		16'b0010101001011100: color_data = 12'b001110100111;
		16'b0010101001011101: color_data = 12'b001110100111;
		16'b0010101001011110: color_data = 12'b001110100111;
		16'b0010101001011111: color_data = 12'b001110100111;
		16'b0010101001100000: color_data = 12'b001110100111;
		16'b0010101001100001: color_data = 12'b001110100111;
		16'b0010101001100010: color_data = 12'b001110100111;
		16'b0010101001100011: color_data = 12'b001110100111;
		16'b0010101001100100: color_data = 12'b001110100111;
		16'b0010101001100101: color_data = 12'b001110100111;
		16'b0010101001100110: color_data = 12'b001110100111;
		16'b0010101001100111: color_data = 12'b001110100111;
		16'b0010101001101000: color_data = 12'b001110100111;
		16'b0010101001101001: color_data = 12'b001110100111;
		16'b0010101001101010: color_data = 12'b001110100111;
		16'b0010101001101011: color_data = 12'b001110100111;
		16'b0010101001101100: color_data = 12'b001110100111;
		16'b0010101001101101: color_data = 12'b001110100111;
		16'b0010101001101110: color_data = 12'b001110100111;
		16'b0010101001110101: color_data = 12'b001110100111;
		16'b0010101001110110: color_data = 12'b001110100111;
		16'b0010101001110111: color_data = 12'b001110100111;
		16'b0010101001111000: color_data = 12'b001110100111;
		16'b0010101001111001: color_data = 12'b001110100111;
		16'b0010101001111010: color_data = 12'b001110100111;
		16'b0010101001111011: color_data = 12'b001110100111;
		16'b0010101001111100: color_data = 12'b001110100111;
		16'b0010101001111101: color_data = 12'b001110100111;
		16'b0010101001111110: color_data = 12'b001110100111;
		16'b0010101001111111: color_data = 12'b001110100111;
		16'b0010101010000000: color_data = 12'b001110100111;
		16'b0010101010000001: color_data = 12'b001110100111;
		16'b0010101010000010: color_data = 12'b001110100111;
		16'b0010101010000011: color_data = 12'b001110100111;
		16'b0010101010000100: color_data = 12'b001110100111;
		16'b0010101010000101: color_data = 12'b001110100111;
		16'b0010101010000110: color_data = 12'b001110100111;
		16'b0010101010000111: color_data = 12'b001110100111;
		16'b0010101010001000: color_data = 12'b001110100111;
		16'b0010101010001001: color_data = 12'b001110100111;
		16'b0010101010001010: color_data = 12'b001110100111;
		16'b0010101010001011: color_data = 12'b001110100111;
		16'b0010101010001100: color_data = 12'b001110100111;
		16'b0010101010001101: color_data = 12'b001110100111;
		16'b0010101010001110: color_data = 12'b001110100111;
		16'b0010101010001111: color_data = 12'b001110100111;
		16'b0010101010010000: color_data = 12'b001110100111;
		16'b0010101010010001: color_data = 12'b001110100111;
		16'b0010101010010010: color_data = 12'b001110100111;
		16'b0010101010010011: color_data = 12'b001110100111;
		16'b0010101010100110: color_data = 12'b001110100111;
		16'b0010101010100111: color_data = 12'b001110100111;
		16'b0010101010101000: color_data = 12'b001110100111;
		16'b0010101010101001: color_data = 12'b001110100111;
		16'b0010101010101010: color_data = 12'b001110100111;
		16'b0010101010101011: color_data = 12'b001110100111;
		16'b0010101010101100: color_data = 12'b001110100111;
		16'b0010101010101101: color_data = 12'b001110100111;
		16'b0010101010101110: color_data = 12'b001110100111;
		16'b0010101010101111: color_data = 12'b001110100111;
		16'b0010101010110000: color_data = 12'b001110100111;
		16'b0010101010110001: color_data = 12'b001110100111;
		16'b0010101010110010: color_data = 12'b001110100111;
		16'b0010101010110011: color_data = 12'b001110100111;
		16'b0010101010110100: color_data = 12'b001110100111;
		16'b0010101010110101: color_data = 12'b001110100111;
		16'b0010101010110110: color_data = 12'b001110100111;
		16'b0010101010110111: color_data = 12'b001110100111;
		16'b0010101010111000: color_data = 12'b001110100111;
		16'b0010101010111001: color_data = 12'b001110100111;
		16'b0010101010111010: color_data = 12'b001110100111;
		16'b0010101010111011: color_data = 12'b001110100111;
		16'b0010101010111100: color_data = 12'b001110100111;
		16'b0010101010111101: color_data = 12'b001110100111;
		16'b0010101010111110: color_data = 12'b001110100111;
		16'b0010101010111111: color_data = 12'b001110100111;
		16'b0010101011000000: color_data = 12'b001110100111;
		16'b0010101011000001: color_data = 12'b001110100111;
		16'b0010101011000010: color_data = 12'b001110100111;
		16'b0010101011000011: color_data = 12'b001110100111;
		16'b0010101011000100: color_data = 12'b001110100111;
		16'b0010101011001011: color_data = 12'b001110100111;
		16'b0010101011001100: color_data = 12'b001110100111;
		16'b0010101011001101: color_data = 12'b001110100111;
		16'b0010101011001110: color_data = 12'b001110100111;
		16'b0010101011001111: color_data = 12'b001110100111;
		16'b0010101011010000: color_data = 12'b001110100111;
		16'b0010101011010001: color_data = 12'b001110100111;
		16'b0010101011010010: color_data = 12'b001110100111;
		16'b0010101011010011: color_data = 12'b001110100111;
		16'b0010101011010100: color_data = 12'b001110100111;
		16'b0010101011010101: color_data = 12'b001110100111;
		16'b0010101011010110: color_data = 12'b001110100111;
		16'b0010101011010111: color_data = 12'b001110100111;
		16'b0010101011011000: color_data = 12'b001110100111;
		16'b0010101011011001: color_data = 12'b001110100111;
		16'b0010101011011010: color_data = 12'b001110100111;
		16'b0010101011011011: color_data = 12'b001110100111;
		16'b0010101011011100: color_data = 12'b001110100111;
		16'b0010101011011101: color_data = 12'b001110100111;
		16'b0010101011011110: color_data = 12'b001110100111;
		16'b0010101011011111: color_data = 12'b001110100111;
		16'b0010101011100000: color_data = 12'b001110100111;
		16'b0010101011100001: color_data = 12'b001110100111;
		16'b0010101011100010: color_data = 12'b001110100111;
		16'b0010101011100011: color_data = 12'b001110100111;
		16'b0010101011100100: color_data = 12'b001110100111;
		16'b0010101011100101: color_data = 12'b001110100111;
		16'b0010101011100110: color_data = 12'b001110100111;
		16'b0010101011100111: color_data = 12'b001110100111;
		16'b0010101011101000: color_data = 12'b001110100111;
		16'b0010101011101001: color_data = 12'b001110100111;
		16'b0010101011101010: color_data = 12'b001110100111;
		16'b0010101011101011: color_data = 12'b001110100111;
		16'b0010101011101100: color_data = 12'b001110100111;
		16'b0010101011101101: color_data = 12'b001110100111;
		16'b0010101011101110: color_data = 12'b001110100111;
		16'b0010101011101111: color_data = 12'b001110100111;
		16'b0010101011110110: color_data = 12'b001110100111;
		16'b0010101011110111: color_data = 12'b001110100111;
		16'b0010101011111000: color_data = 12'b001110100111;
		16'b0010101011111001: color_data = 12'b001110100111;
		16'b0010101011111010: color_data = 12'b001110100111;
		16'b0010101011111011: color_data = 12'b001110100111;
		16'b0010101011111100: color_data = 12'b001110100111;
		16'b0010101011111101: color_data = 12'b001110100111;
		16'b0010101011111110: color_data = 12'b001110100111;
		16'b0010101011111111: color_data = 12'b001110100111;
		16'b0010101100000000: color_data = 12'b001110100111;
		16'b0010101100000001: color_data = 12'b001110100111;
		16'b0010101100000010: color_data = 12'b001110100111;
		16'b0010101100000011: color_data = 12'b001110100111;
		16'b0010101100000100: color_data = 12'b001110100111;
		16'b0010101100000101: color_data = 12'b001110100111;
		16'b0010101100000110: color_data = 12'b001110100111;
		16'b0010101100000111: color_data = 12'b001110100111;
		16'b0010101100001000: color_data = 12'b001110100111;
		16'b0010101100001001: color_data = 12'b001110100111;
		16'b0010101100001010: color_data = 12'b001110100111;
		16'b0010101100001011: color_data = 12'b001110100111;
		16'b0010101100001100: color_data = 12'b001110100111;
		16'b0010101100001101: color_data = 12'b001110100111;
		16'b0010101100001110: color_data = 12'b001110100111;
		16'b0010101100001111: color_data = 12'b001110100111;
		16'b0010101100010000: color_data = 12'b001110100111;
		16'b0010101100010001: color_data = 12'b001110100111;
		16'b0010101100010010: color_data = 12'b001110100111;
		16'b0010101100010011: color_data = 12'b001110100111;
		16'b0010101100010100: color_data = 12'b001110100111;
		16'b0010101100010101: color_data = 12'b001110100111;
		16'b0010101100010110: color_data = 12'b001110100111;
		16'b0010101100010111: color_data = 12'b001110100111;
		16'b0010101100011000: color_data = 12'b001110100111;
		16'b0010101100011001: color_data = 12'b001110100111;
		16'b0010101100011010: color_data = 12'b001110100111;
		16'b0010101100011011: color_data = 12'b001110100111;
		16'b0010101100011100: color_data = 12'b001110100111;
		16'b0010101100011101: color_data = 12'b001110100111;
		16'b0010101100011110: color_data = 12'b001110100111;
		16'b0010101100011111: color_data = 12'b001110100111;
		16'b0010101100100000: color_data = 12'b001110100111;
		16'b0010101100100001: color_data = 12'b001110100111;
		16'b0010101100100010: color_data = 12'b001110100111;
		16'b0010101100100011: color_data = 12'b001110100111;
		16'b0010101100100100: color_data = 12'b001110100111;
		16'b0010101100100101: color_data = 12'b001110100111;
		16'b0010101100100110: color_data = 12'b001110100111;
		16'b0010101100101101: color_data = 12'b001110100111;
		16'b0010101100101110: color_data = 12'b001110100111;
		16'b0010101100101111: color_data = 12'b001110100111;
		16'b0010101100110000: color_data = 12'b001110100111;
		16'b0010101100110001: color_data = 12'b001110100111;
		16'b0010101100110010: color_data = 12'b001110100111;
		16'b0010101100110011: color_data = 12'b001110100111;
		16'b0010101100110100: color_data = 12'b001110100111;
		16'b0010101100110101: color_data = 12'b001110100111;
		16'b0010101100110110: color_data = 12'b001110100111;
		16'b0010101100110111: color_data = 12'b001110100111;
		16'b0010101100111000: color_data = 12'b001110100111;
		16'b0010101100111001: color_data = 12'b001110100111;
		16'b0010101100111010: color_data = 12'b001110100111;
		16'b0010101100111011: color_data = 12'b001110100111;
		16'b0010101100111100: color_data = 12'b001110100111;
		16'b0010101100111101: color_data = 12'b001110100111;
		16'b0010101100111110: color_data = 12'b001110100111;
		16'b0010101100111111: color_data = 12'b001110100111;
		16'b0010101101000000: color_data = 12'b001110100111;
		16'b0010101101000001: color_data = 12'b001110100111;
		16'b0010101101000010: color_data = 12'b001110100111;
		16'b0010101101000011: color_data = 12'b001110100111;
		16'b0010101101000100: color_data = 12'b001110100111;
		16'b0010101101000101: color_data = 12'b001110100111;
		16'b0010101101000110: color_data = 12'b001110100111;
		16'b0010101101000111: color_data = 12'b001110100111;
		16'b0010101101001000: color_data = 12'b001110100111;
		16'b0010101101001001: color_data = 12'b001110100111;
		16'b0010101101001010: color_data = 12'b001110100111;
		16'b0010101101011110: color_data = 12'b001110100111;
		16'b0010101101011111: color_data = 12'b001110100111;
		16'b0010101101100000: color_data = 12'b001110100111;
		16'b0010101101100001: color_data = 12'b001110100111;
		16'b0010101101100010: color_data = 12'b001110100111;
		16'b0010101101100011: color_data = 12'b001110100111;
		16'b0010101101100100: color_data = 12'b001110100111;
		16'b0010101101100101: color_data = 12'b001110100111;
		16'b0010101101100110: color_data = 12'b001110100111;
		16'b0010101101100111: color_data = 12'b001110100111;
		16'b0010101101101000: color_data = 12'b001110100111;
		16'b0010101101101001: color_data = 12'b001110100111;
		16'b0010101101101010: color_data = 12'b001110100111;
		16'b0010101101101011: color_data = 12'b001110100111;
		16'b0010101101101100: color_data = 12'b001110100111;
		16'b0010101101101101: color_data = 12'b001110100111;
		16'b0010101101101110: color_data = 12'b001110100111;
		16'b0010101101101111: color_data = 12'b001110100111;
		16'b0010101101110000: color_data = 12'b001110100111;
		16'b0010101101110001: color_data = 12'b001110100111;
		16'b0010101101110010: color_data = 12'b001110100111;
		16'b0010101101110011: color_data = 12'b001110100111;
		16'b0010101101110100: color_data = 12'b001110100111;
		16'b0010101101110101: color_data = 12'b001110100111;
		16'b0010101101110110: color_data = 12'b001110100111;
		16'b0010101101110111: color_data = 12'b001110100111;
		16'b0010101101111000: color_data = 12'b001110100111;
		16'b0010101101111001: color_data = 12'b001110100111;
		16'b0010101101111010: color_data = 12'b001110100111;
		16'b0010101101111011: color_data = 12'b001110100111;
		16'b0010110000000111: color_data = 12'b001110100111;
		16'b0010110000001000: color_data = 12'b001110100111;
		16'b0010110000001001: color_data = 12'b001110100111;
		16'b0010110000001010: color_data = 12'b001110100111;
		16'b0010110000001011: color_data = 12'b001110100111;
		16'b0010110000001100: color_data = 12'b001110100111;
		16'b0010110000001101: color_data = 12'b001110100111;
		16'b0010110000001110: color_data = 12'b001110100111;
		16'b0010110000001111: color_data = 12'b001110100111;
		16'b0010110000010000: color_data = 12'b001110100111;
		16'b0010110000010001: color_data = 12'b001110100111;
		16'b0010110000010010: color_data = 12'b001110100111;
		16'b0010110000010011: color_data = 12'b001110100111;
		16'b0010110000010100: color_data = 12'b001110100111;
		16'b0010110000010101: color_data = 12'b001110100111;
		16'b0010110000010110: color_data = 12'b001110100111;
		16'b0010110000010111: color_data = 12'b001110100111;
		16'b0010110000011000: color_data = 12'b001110100111;
		16'b0010110000011001: color_data = 12'b001110100111;
		16'b0010110000011010: color_data = 12'b001110100111;
		16'b0010110000011011: color_data = 12'b001110100111;
		16'b0010110000011100: color_data = 12'b001110100111;
		16'b0010110000011101: color_data = 12'b001110100111;
		16'b0010110000011110: color_data = 12'b001110100111;
		16'b0010110000011111: color_data = 12'b001110100111;
		16'b0010110000100000: color_data = 12'b001110100111;
		16'b0010110000100001: color_data = 12'b001110100111;
		16'b0010110000100010: color_data = 12'b001110100111;
		16'b0010110000100011: color_data = 12'b001110100111;
		16'b0010110000100100: color_data = 12'b001110100111;
		16'b0010110000101011: color_data = 12'b001110100111;
		16'b0010110000101100: color_data = 12'b001110100111;
		16'b0010110000101101: color_data = 12'b001110100111;
		16'b0010110000101110: color_data = 12'b001110100111;
		16'b0010110000101111: color_data = 12'b001110100111;
		16'b0010110000110000: color_data = 12'b001110100111;
		16'b0010110000110001: color_data = 12'b001110100111;
		16'b0010110000110010: color_data = 12'b001110100111;
		16'b0010110000110011: color_data = 12'b001110100111;
		16'b0010110000110100: color_data = 12'b001110100111;
		16'b0010110000110101: color_data = 12'b001110100111;
		16'b0010110000110110: color_data = 12'b001110100111;
		16'b0010110000110111: color_data = 12'b001110100111;
		16'b0010110001000100: color_data = 12'b001110100111;
		16'b0010110001000101: color_data = 12'b001110100111;
		16'b0010110001000110: color_data = 12'b001110100111;
		16'b0010110001000111: color_data = 12'b001110100111;
		16'b0010110001001000: color_data = 12'b001110100111;
		16'b0010110001001001: color_data = 12'b001110100111;
		16'b0010110001001010: color_data = 12'b001110100111;
		16'b0010110001001011: color_data = 12'b001110100111;
		16'b0010110001001100: color_data = 12'b001110100111;
		16'b0010110001001101: color_data = 12'b001110100111;
		16'b0010110001001110: color_data = 12'b001110100111;
		16'b0010110001001111: color_data = 12'b001110100111;
		16'b0010110001010110: color_data = 12'b001110100111;
		16'b0010110001010111: color_data = 12'b001110100111;
		16'b0010110001011000: color_data = 12'b001110100111;
		16'b0010110001011001: color_data = 12'b001110100111;
		16'b0010110001011010: color_data = 12'b001110100111;
		16'b0010110001011011: color_data = 12'b001110100111;
		16'b0010110001011100: color_data = 12'b001110100111;
		16'b0010110001011101: color_data = 12'b001110100111;
		16'b0010110001011110: color_data = 12'b001110100111;
		16'b0010110001011111: color_data = 12'b001110100111;
		16'b0010110001100000: color_data = 12'b001110100111;
		16'b0010110001100001: color_data = 12'b001110100111;
		16'b0010110001100010: color_data = 12'b001110100111;
		16'b0010110001100011: color_data = 12'b001110100111;
		16'b0010110001100100: color_data = 12'b001110100111;
		16'b0010110001100101: color_data = 12'b001110100111;
		16'b0010110001100110: color_data = 12'b001110100111;
		16'b0010110001100111: color_data = 12'b001110100111;
		16'b0010110001101000: color_data = 12'b001110100111;
		16'b0010110001101001: color_data = 12'b001110100111;
		16'b0010110001101010: color_data = 12'b001110100111;
		16'b0010110001101011: color_data = 12'b001110100111;
		16'b0010110001101100: color_data = 12'b001110100111;
		16'b0010110001101101: color_data = 12'b001110100111;
		16'b0010110001101110: color_data = 12'b001110100111;
		16'b0010110001110101: color_data = 12'b001110100111;
		16'b0010110001110110: color_data = 12'b001110100111;
		16'b0010110001110111: color_data = 12'b001110100111;
		16'b0010110001111000: color_data = 12'b001110100111;
		16'b0010110001111001: color_data = 12'b001110100111;
		16'b0010110001111010: color_data = 12'b001110100111;
		16'b0010110001111011: color_data = 12'b001110100111;
		16'b0010110001111100: color_data = 12'b001110100111;
		16'b0010110001111101: color_data = 12'b001110100111;
		16'b0010110001111110: color_data = 12'b001110100111;
		16'b0010110001111111: color_data = 12'b001110100111;
		16'b0010110010000000: color_data = 12'b001110100111;
		16'b0010110010000001: color_data = 12'b001110100111;
		16'b0010110010000010: color_data = 12'b001110100111;
		16'b0010110010000011: color_data = 12'b001110100111;
		16'b0010110010000100: color_data = 12'b001110100111;
		16'b0010110010000101: color_data = 12'b001110100111;
		16'b0010110010000110: color_data = 12'b001110100111;
		16'b0010110010000111: color_data = 12'b001110100111;
		16'b0010110010001000: color_data = 12'b001110100111;
		16'b0010110010001001: color_data = 12'b001110100111;
		16'b0010110010001010: color_data = 12'b001110100111;
		16'b0010110010001011: color_data = 12'b001110100111;
		16'b0010110010001100: color_data = 12'b001110100111;
		16'b0010110010001101: color_data = 12'b001110100111;
		16'b0010110010001110: color_data = 12'b001110100111;
		16'b0010110010001111: color_data = 12'b001110100111;
		16'b0010110010010000: color_data = 12'b001110100111;
		16'b0010110010010001: color_data = 12'b001110100111;
		16'b0010110010010010: color_data = 12'b001110100111;
		16'b0010110010010011: color_data = 12'b001110100111;
		16'b0010110010100110: color_data = 12'b001110100111;
		16'b0010110010100111: color_data = 12'b001110100111;
		16'b0010110010101000: color_data = 12'b001110100111;
		16'b0010110010101001: color_data = 12'b001110100111;
		16'b0010110010101010: color_data = 12'b001110100111;
		16'b0010110010101011: color_data = 12'b001110100111;
		16'b0010110010101100: color_data = 12'b001110100111;
		16'b0010110010101101: color_data = 12'b001110100111;
		16'b0010110010101110: color_data = 12'b001110100111;
		16'b0010110010101111: color_data = 12'b001110100111;
		16'b0010110010110000: color_data = 12'b001110100111;
		16'b0010110010110001: color_data = 12'b001110100111;
		16'b0010110010110010: color_data = 12'b001110100111;
		16'b0010110010110011: color_data = 12'b001110100111;
		16'b0010110010110100: color_data = 12'b001110100111;
		16'b0010110010110101: color_data = 12'b001110100111;
		16'b0010110010110110: color_data = 12'b001110100111;
		16'b0010110010110111: color_data = 12'b001110100111;
		16'b0010110010111000: color_data = 12'b001110100111;
		16'b0010110010111001: color_data = 12'b001110100111;
		16'b0010110010111010: color_data = 12'b001110100111;
		16'b0010110010111011: color_data = 12'b001110100111;
		16'b0010110010111100: color_data = 12'b001110100111;
		16'b0010110010111101: color_data = 12'b001110100111;
		16'b0010110010111110: color_data = 12'b001110100111;
		16'b0010110010111111: color_data = 12'b001110100111;
		16'b0010110011000000: color_data = 12'b001110100111;
		16'b0010110011000001: color_data = 12'b001110100111;
		16'b0010110011000010: color_data = 12'b001110100111;
		16'b0010110011000011: color_data = 12'b001110100111;
		16'b0010110011000100: color_data = 12'b001110100111;
		16'b0010110011001011: color_data = 12'b001110100111;
		16'b0010110011001100: color_data = 12'b001110100111;
		16'b0010110011001101: color_data = 12'b001110100111;
		16'b0010110011001110: color_data = 12'b001110100111;
		16'b0010110011001111: color_data = 12'b001110100111;
		16'b0010110011010000: color_data = 12'b001110100111;
		16'b0010110011010001: color_data = 12'b001110100111;
		16'b0010110011010010: color_data = 12'b001110100111;
		16'b0010110011010011: color_data = 12'b001110100111;
		16'b0010110011010100: color_data = 12'b001110100111;
		16'b0010110011010101: color_data = 12'b001110100111;
		16'b0010110011010110: color_data = 12'b001110100111;
		16'b0010110011010111: color_data = 12'b001110100111;
		16'b0010110011011000: color_data = 12'b001110100111;
		16'b0010110011011001: color_data = 12'b001110100111;
		16'b0010110011011010: color_data = 12'b001110100111;
		16'b0010110011011011: color_data = 12'b001110100111;
		16'b0010110011011100: color_data = 12'b001110100111;
		16'b0010110011011101: color_data = 12'b001110100111;
		16'b0010110011011110: color_data = 12'b001110100111;
		16'b0010110011011111: color_data = 12'b001110100111;
		16'b0010110011100000: color_data = 12'b001110100111;
		16'b0010110011100001: color_data = 12'b001110100111;
		16'b0010110011100010: color_data = 12'b001110100111;
		16'b0010110011100011: color_data = 12'b001110100111;
		16'b0010110011100100: color_data = 12'b001110100111;
		16'b0010110011100101: color_data = 12'b001110100111;
		16'b0010110011100110: color_data = 12'b001110100111;
		16'b0010110011100111: color_data = 12'b001110100111;
		16'b0010110011101000: color_data = 12'b001110100111;
		16'b0010110011101001: color_data = 12'b001110100111;
		16'b0010110011101010: color_data = 12'b001110100111;
		16'b0010110011101011: color_data = 12'b001110100111;
		16'b0010110011101100: color_data = 12'b001110100111;
		16'b0010110011101101: color_data = 12'b001110100111;
		16'b0010110011101110: color_data = 12'b001110100111;
		16'b0010110011101111: color_data = 12'b001110100111;
		16'b0010110011110110: color_data = 12'b001110100111;
		16'b0010110011110111: color_data = 12'b001110100111;
		16'b0010110011111000: color_data = 12'b001110100111;
		16'b0010110011111001: color_data = 12'b001110100111;
		16'b0010110011111010: color_data = 12'b001110100111;
		16'b0010110011111011: color_data = 12'b001110100111;
		16'b0010110011111100: color_data = 12'b001110100111;
		16'b0010110011111101: color_data = 12'b001110100111;
		16'b0010110011111110: color_data = 12'b001110100111;
		16'b0010110011111111: color_data = 12'b001110100111;
		16'b0010110100000000: color_data = 12'b001110100111;
		16'b0010110100000001: color_data = 12'b001110100111;
		16'b0010110100000010: color_data = 12'b001110100111;
		16'b0010110100000011: color_data = 12'b001110100111;
		16'b0010110100000100: color_data = 12'b001110100111;
		16'b0010110100000101: color_data = 12'b001110100111;
		16'b0010110100000110: color_data = 12'b001110100111;
		16'b0010110100000111: color_data = 12'b001110100111;
		16'b0010110100001000: color_data = 12'b001110100111;
		16'b0010110100001001: color_data = 12'b001110100111;
		16'b0010110100001010: color_data = 12'b001110100111;
		16'b0010110100001011: color_data = 12'b001110100111;
		16'b0010110100001100: color_data = 12'b001110100111;
		16'b0010110100001101: color_data = 12'b001110100111;
		16'b0010110100001110: color_data = 12'b001110100111;
		16'b0010110100001111: color_data = 12'b001110100111;
		16'b0010110100010000: color_data = 12'b001110100111;
		16'b0010110100010001: color_data = 12'b001110100111;
		16'b0010110100010010: color_data = 12'b001110100111;
		16'b0010110100010011: color_data = 12'b001110100111;
		16'b0010110100010100: color_data = 12'b001110100111;
		16'b0010110100010101: color_data = 12'b001110100111;
		16'b0010110100010110: color_data = 12'b001110100111;
		16'b0010110100010111: color_data = 12'b001110100111;
		16'b0010110100011000: color_data = 12'b001110100111;
		16'b0010110100011001: color_data = 12'b001110100111;
		16'b0010110100011010: color_data = 12'b001110100111;
		16'b0010110100011011: color_data = 12'b001110100111;
		16'b0010110100011100: color_data = 12'b001110100111;
		16'b0010110100011101: color_data = 12'b001110100111;
		16'b0010110100011110: color_data = 12'b001110100111;
		16'b0010110100011111: color_data = 12'b001110100111;
		16'b0010110100100000: color_data = 12'b001110100111;
		16'b0010110100100001: color_data = 12'b001110100111;
		16'b0010110100100010: color_data = 12'b001110100111;
		16'b0010110100100011: color_data = 12'b001110100111;
		16'b0010110100100100: color_data = 12'b001110100111;
		16'b0010110100100101: color_data = 12'b001110100111;
		16'b0010110100100110: color_data = 12'b001110100111;
		16'b0010110100101101: color_data = 12'b001110100111;
		16'b0010110100101110: color_data = 12'b001110100111;
		16'b0010110100101111: color_data = 12'b001110100111;
		16'b0010110100110000: color_data = 12'b001110100111;
		16'b0010110100110001: color_data = 12'b001110100111;
		16'b0010110100110010: color_data = 12'b001110100111;
		16'b0010110100110011: color_data = 12'b001110100111;
		16'b0010110100110100: color_data = 12'b001110100111;
		16'b0010110100110101: color_data = 12'b001110100111;
		16'b0010110100110110: color_data = 12'b001110100111;
		16'b0010110100110111: color_data = 12'b001110100111;
		16'b0010110100111000: color_data = 12'b001110100111;
		16'b0010110100111001: color_data = 12'b001110100111;
		16'b0010110100111010: color_data = 12'b001110100111;
		16'b0010110100111011: color_data = 12'b001110100111;
		16'b0010110100111100: color_data = 12'b001110100111;
		16'b0010110100111101: color_data = 12'b001110100111;
		16'b0010110100111110: color_data = 12'b001110100111;
		16'b0010110100111111: color_data = 12'b001110100111;
		16'b0010110101000000: color_data = 12'b001110100111;
		16'b0010110101000001: color_data = 12'b001110100111;
		16'b0010110101000010: color_data = 12'b001110100111;
		16'b0010110101000011: color_data = 12'b001110100111;
		16'b0010110101000100: color_data = 12'b001110100111;
		16'b0010110101000101: color_data = 12'b001110100111;
		16'b0010110101000110: color_data = 12'b001110100111;
		16'b0010110101000111: color_data = 12'b001110100111;
		16'b0010110101001000: color_data = 12'b001110100111;
		16'b0010110101001001: color_data = 12'b001110100111;
		16'b0010110101001010: color_data = 12'b001110100111;
		16'b0010110101011110: color_data = 12'b001110100111;
		16'b0010110101011111: color_data = 12'b001110100111;
		16'b0010110101100000: color_data = 12'b001110100111;
		16'b0010110101100001: color_data = 12'b001110100111;
		16'b0010110101100010: color_data = 12'b001110100111;
		16'b0010110101100011: color_data = 12'b001110100111;
		16'b0010110101100100: color_data = 12'b001110100111;
		16'b0010110101100101: color_data = 12'b001110100111;
		16'b0010110101100110: color_data = 12'b001110100111;
		16'b0010110101100111: color_data = 12'b001110100111;
		16'b0010110101101000: color_data = 12'b001110100111;
		16'b0010110101101001: color_data = 12'b001110100111;
		16'b0010110101101010: color_data = 12'b001110100111;
		16'b0010110101101011: color_data = 12'b001110100111;
		16'b0010110101101100: color_data = 12'b001110100111;
		16'b0010110101101101: color_data = 12'b001110100111;
		16'b0010110101101110: color_data = 12'b001110100111;
		16'b0010110101101111: color_data = 12'b001110100111;
		16'b0010110101110000: color_data = 12'b001110100111;
		16'b0010110101110001: color_data = 12'b001110100111;
		16'b0010110101110010: color_data = 12'b001110100111;
		16'b0010110101110011: color_data = 12'b001110100111;
		16'b0010110101110100: color_data = 12'b001110100111;
		16'b0010110101110101: color_data = 12'b001110100111;
		16'b0010110101110110: color_data = 12'b001110100111;
		16'b0010110101110111: color_data = 12'b001110100111;
		16'b0010110101111000: color_data = 12'b001110100111;
		16'b0010110101111001: color_data = 12'b001110100111;
		16'b0010110101111010: color_data = 12'b001110100111;
		16'b0010110101111011: color_data = 12'b001110100111;
		16'b0010111000000111: color_data = 12'b001110100111;
		16'b0010111000001000: color_data = 12'b001110100111;
		16'b0010111000001001: color_data = 12'b001110100111;
		16'b0010111000001010: color_data = 12'b001110100111;
		16'b0010111000001011: color_data = 12'b001110100111;
		16'b0010111000001100: color_data = 12'b001110100111;
		16'b0010111000001101: color_data = 12'b001110100111;
		16'b0010111000001110: color_data = 12'b001110100111;
		16'b0010111000001111: color_data = 12'b001110100111;
		16'b0010111000010000: color_data = 12'b001110100111;
		16'b0010111000010001: color_data = 12'b001110100111;
		16'b0010111000010010: color_data = 12'b001110100111;
		16'b0010111000010011: color_data = 12'b001110100111;
		16'b0010111000010100: color_data = 12'b001110100111;
		16'b0010111000010101: color_data = 12'b001110100111;
		16'b0010111000010110: color_data = 12'b001110100111;
		16'b0010111000010111: color_data = 12'b001110100111;
		16'b0010111000011000: color_data = 12'b001110100111;
		16'b0010111000011001: color_data = 12'b001110100111;
		16'b0010111000011010: color_data = 12'b001110100111;
		16'b0010111000011011: color_data = 12'b001110100111;
		16'b0010111000011100: color_data = 12'b001110100111;
		16'b0010111000011101: color_data = 12'b001110100111;
		16'b0010111000011110: color_data = 12'b001110100111;
		16'b0010111000011111: color_data = 12'b001110100111;
		16'b0010111000100000: color_data = 12'b001110100111;
		16'b0010111000100001: color_data = 12'b001110100111;
		16'b0010111000100010: color_data = 12'b001110100111;
		16'b0010111000100011: color_data = 12'b001110100111;
		16'b0010111000100100: color_data = 12'b001110100111;
		16'b0010111000101011: color_data = 12'b001110100111;
		16'b0010111000101100: color_data = 12'b001110100111;
		16'b0010111000101101: color_data = 12'b001110100111;
		16'b0010111000101110: color_data = 12'b001110100111;
		16'b0010111000101111: color_data = 12'b001110100111;
		16'b0010111000110000: color_data = 12'b001110100111;
		16'b0010111000110001: color_data = 12'b001110100111;
		16'b0010111000110010: color_data = 12'b001110100111;
		16'b0010111000110011: color_data = 12'b001110100111;
		16'b0010111000110100: color_data = 12'b001110100111;
		16'b0010111000110101: color_data = 12'b001110100111;
		16'b0010111000110110: color_data = 12'b001110100111;
		16'b0010111000110111: color_data = 12'b001110100111;
		16'b0010111001000100: color_data = 12'b001110100111;
		16'b0010111001000101: color_data = 12'b001110100111;
		16'b0010111001000110: color_data = 12'b001110100111;
		16'b0010111001000111: color_data = 12'b001110100111;
		16'b0010111001001000: color_data = 12'b001110100111;
		16'b0010111001001001: color_data = 12'b001110100111;
		16'b0010111001001010: color_data = 12'b001110100111;
		16'b0010111001001011: color_data = 12'b001110100111;
		16'b0010111001001100: color_data = 12'b001110100111;
		16'b0010111001001101: color_data = 12'b001110100111;
		16'b0010111001001110: color_data = 12'b001110100111;
		16'b0010111001001111: color_data = 12'b001110100111;
		16'b0010111001010110: color_data = 12'b001110100111;
		16'b0010111001010111: color_data = 12'b001110100111;
		16'b0010111001011000: color_data = 12'b001110100111;
		16'b0010111001011001: color_data = 12'b001110100111;
		16'b0010111001011010: color_data = 12'b001110100111;
		16'b0010111001011011: color_data = 12'b001110100111;
		16'b0010111001011100: color_data = 12'b001110100111;
		16'b0010111001011101: color_data = 12'b001110100111;
		16'b0010111001011110: color_data = 12'b001110100111;
		16'b0010111001011111: color_data = 12'b001110100111;
		16'b0010111001100000: color_data = 12'b001110100111;
		16'b0010111001100001: color_data = 12'b001110100111;
		16'b0010111001100010: color_data = 12'b001110100111;
		16'b0010111001100011: color_data = 12'b001110100111;
		16'b0010111001100100: color_data = 12'b001110100111;
		16'b0010111001100101: color_data = 12'b001110100111;
		16'b0010111001100110: color_data = 12'b001110100111;
		16'b0010111001100111: color_data = 12'b001110100111;
		16'b0010111001101000: color_data = 12'b001110100111;
		16'b0010111001101001: color_data = 12'b001110100111;
		16'b0010111001101010: color_data = 12'b001110100111;
		16'b0010111001101011: color_data = 12'b001110100111;
		16'b0010111001101100: color_data = 12'b001110100111;
		16'b0010111001101101: color_data = 12'b001110100111;
		16'b0010111001101110: color_data = 12'b001110100111;
		16'b0010111001110101: color_data = 12'b001110100111;
		16'b0010111001110110: color_data = 12'b001110100111;
		16'b0010111001110111: color_data = 12'b001110100111;
		16'b0010111001111000: color_data = 12'b001110100111;
		16'b0010111001111001: color_data = 12'b001110100111;
		16'b0010111001111010: color_data = 12'b001110100111;
		16'b0010111001111011: color_data = 12'b001110100111;
		16'b0010111001111100: color_data = 12'b001110100111;
		16'b0010111001111101: color_data = 12'b001110100111;
		16'b0010111001111110: color_data = 12'b001110100111;
		16'b0010111001111111: color_data = 12'b001110100111;
		16'b0010111010000000: color_data = 12'b001110100111;
		16'b0010111010000001: color_data = 12'b001110100111;
		16'b0010111010000010: color_data = 12'b001110100111;
		16'b0010111010000011: color_data = 12'b001110100111;
		16'b0010111010000100: color_data = 12'b001110100111;
		16'b0010111010000101: color_data = 12'b001110100111;
		16'b0010111010000110: color_data = 12'b001110100111;
		16'b0010111010000111: color_data = 12'b001110100111;
		16'b0010111010001000: color_data = 12'b001110100111;
		16'b0010111010001001: color_data = 12'b001110100111;
		16'b0010111010001010: color_data = 12'b001110100111;
		16'b0010111010001011: color_data = 12'b001110100111;
		16'b0010111010001100: color_data = 12'b001110100111;
		16'b0010111010001101: color_data = 12'b001110100111;
		16'b0010111010001110: color_data = 12'b001110100111;
		16'b0010111010001111: color_data = 12'b001110100111;
		16'b0010111010010000: color_data = 12'b001110100111;
		16'b0010111010010001: color_data = 12'b001110100111;
		16'b0010111010010010: color_data = 12'b001110100111;
		16'b0010111010010011: color_data = 12'b001110100111;
		16'b0010111010100110: color_data = 12'b001110100111;
		16'b0010111010100111: color_data = 12'b001110100111;
		16'b0010111010101000: color_data = 12'b001110100111;
		16'b0010111010101001: color_data = 12'b001110100111;
		16'b0010111010101010: color_data = 12'b001110100111;
		16'b0010111010101011: color_data = 12'b001110100111;
		16'b0010111010101100: color_data = 12'b001110100111;
		16'b0010111010101101: color_data = 12'b001110100111;
		16'b0010111010101110: color_data = 12'b001110100111;
		16'b0010111010101111: color_data = 12'b001110100111;
		16'b0010111010110000: color_data = 12'b001110100111;
		16'b0010111010110001: color_data = 12'b001110100111;
		16'b0010111010110010: color_data = 12'b001110100111;
		16'b0010111010110011: color_data = 12'b001110100111;
		16'b0010111010110100: color_data = 12'b001110100111;
		16'b0010111010110101: color_data = 12'b001110100111;
		16'b0010111010110110: color_data = 12'b001110100111;
		16'b0010111010110111: color_data = 12'b001110100111;
		16'b0010111010111000: color_data = 12'b001110100111;
		16'b0010111010111001: color_data = 12'b001110100111;
		16'b0010111010111010: color_data = 12'b001110100111;
		16'b0010111010111011: color_data = 12'b001110100111;
		16'b0010111010111100: color_data = 12'b001110100111;
		16'b0010111010111101: color_data = 12'b001110100111;
		16'b0010111010111110: color_data = 12'b001110100111;
		16'b0010111010111111: color_data = 12'b001110100111;
		16'b0010111011000000: color_data = 12'b001110100111;
		16'b0010111011000001: color_data = 12'b001110100111;
		16'b0010111011000010: color_data = 12'b001110100111;
		16'b0010111011000011: color_data = 12'b001110100111;
		16'b0010111011000100: color_data = 12'b001110100111;
		16'b0010111011001011: color_data = 12'b001110100111;
		16'b0010111011001100: color_data = 12'b001110100111;
		16'b0010111011001101: color_data = 12'b001110100111;
		16'b0010111011001110: color_data = 12'b001110100111;
		16'b0010111011001111: color_data = 12'b001110100111;
		16'b0010111011010000: color_data = 12'b001110100111;
		16'b0010111011010001: color_data = 12'b001110100111;
		16'b0010111011010010: color_data = 12'b001110100111;
		16'b0010111011010011: color_data = 12'b001110100111;
		16'b0010111011010100: color_data = 12'b001110100111;
		16'b0010111011010101: color_data = 12'b001110100111;
		16'b0010111011010110: color_data = 12'b001110100111;
		16'b0010111011010111: color_data = 12'b001110100111;
		16'b0010111011011000: color_data = 12'b001110100111;
		16'b0010111011011001: color_data = 12'b001110100111;
		16'b0010111011011010: color_data = 12'b001110100111;
		16'b0010111011011011: color_data = 12'b001110100111;
		16'b0010111011011100: color_data = 12'b001110100111;
		16'b0010111011011101: color_data = 12'b001110100111;
		16'b0010111011011110: color_data = 12'b001110100111;
		16'b0010111011011111: color_data = 12'b001110100111;
		16'b0010111011100000: color_data = 12'b001110100111;
		16'b0010111011100001: color_data = 12'b001110100111;
		16'b0010111011100010: color_data = 12'b001110100111;
		16'b0010111011100011: color_data = 12'b001110100111;
		16'b0010111011100100: color_data = 12'b001110100111;
		16'b0010111011100101: color_data = 12'b001110100111;
		16'b0010111011100110: color_data = 12'b001110100111;
		16'b0010111011100111: color_data = 12'b001110100111;
		16'b0010111011101000: color_data = 12'b001110100111;
		16'b0010111011101001: color_data = 12'b001110100111;
		16'b0010111011101010: color_data = 12'b001110100111;
		16'b0010111011101011: color_data = 12'b001110100111;
		16'b0010111011101100: color_data = 12'b001110100111;
		16'b0010111011101101: color_data = 12'b001110100111;
		16'b0010111011101110: color_data = 12'b001110100111;
		16'b0010111011101111: color_data = 12'b001110100111;
		16'b0010111011110110: color_data = 12'b001110100111;
		16'b0010111011110111: color_data = 12'b001110100111;
		16'b0010111011111000: color_data = 12'b001110100111;
		16'b0010111011111001: color_data = 12'b001110100111;
		16'b0010111011111010: color_data = 12'b001110100111;
		16'b0010111011111011: color_data = 12'b001110100111;
		16'b0010111011111100: color_data = 12'b001110100111;
		16'b0010111011111101: color_data = 12'b001110100111;
		16'b0010111011111110: color_data = 12'b001110100111;
		16'b0010111011111111: color_data = 12'b001110100111;
		16'b0010111100000000: color_data = 12'b001110100111;
		16'b0010111100000001: color_data = 12'b001110100111;
		16'b0010111100000010: color_data = 12'b001110100111;
		16'b0010111100000011: color_data = 12'b001110100111;
		16'b0010111100000100: color_data = 12'b001110100111;
		16'b0010111100000101: color_data = 12'b001110100111;
		16'b0010111100000110: color_data = 12'b001110100111;
		16'b0010111100000111: color_data = 12'b001110100111;
		16'b0010111100001000: color_data = 12'b001110100111;
		16'b0010111100001001: color_data = 12'b001110100111;
		16'b0010111100001010: color_data = 12'b001110100111;
		16'b0010111100001011: color_data = 12'b001110100111;
		16'b0010111100001100: color_data = 12'b001110100111;
		16'b0010111100001101: color_data = 12'b001110100111;
		16'b0010111100001110: color_data = 12'b001110100111;
		16'b0010111100001111: color_data = 12'b001110100111;
		16'b0010111100010000: color_data = 12'b001110100111;
		16'b0010111100010001: color_data = 12'b001110100111;
		16'b0010111100010010: color_data = 12'b001110100111;
		16'b0010111100010011: color_data = 12'b001110100111;
		16'b0010111100010100: color_data = 12'b001110100111;
		16'b0010111100010101: color_data = 12'b001110100111;
		16'b0010111100010110: color_data = 12'b001110100111;
		16'b0010111100010111: color_data = 12'b001110100111;
		16'b0010111100011000: color_data = 12'b001110100111;
		16'b0010111100011001: color_data = 12'b001110100111;
		16'b0010111100011010: color_data = 12'b001110100111;
		16'b0010111100011011: color_data = 12'b001110100111;
		16'b0010111100011100: color_data = 12'b001110100111;
		16'b0010111100011101: color_data = 12'b001110100111;
		16'b0010111100011110: color_data = 12'b001110100111;
		16'b0010111100011111: color_data = 12'b001110100111;
		16'b0010111100100000: color_data = 12'b001110100111;
		16'b0010111100100001: color_data = 12'b001110100111;
		16'b0010111100100010: color_data = 12'b001110100111;
		16'b0010111100100011: color_data = 12'b001110100111;
		16'b0010111100100100: color_data = 12'b001110100111;
		16'b0010111100100101: color_data = 12'b001110100111;
		16'b0010111100100110: color_data = 12'b001110100111;
		16'b0010111100101101: color_data = 12'b001110100111;
		16'b0010111100101110: color_data = 12'b001110100111;
		16'b0010111100101111: color_data = 12'b001110100111;
		16'b0010111100110000: color_data = 12'b001110100111;
		16'b0010111100110001: color_data = 12'b001110100111;
		16'b0010111100110010: color_data = 12'b001110100111;
		16'b0010111100110011: color_data = 12'b001110100111;
		16'b0010111100110100: color_data = 12'b001110100111;
		16'b0010111100110101: color_data = 12'b001110100111;
		16'b0010111100110110: color_data = 12'b001110100111;
		16'b0010111100110111: color_data = 12'b001110100111;
		16'b0010111100111000: color_data = 12'b001110100111;
		16'b0010111100111001: color_data = 12'b001110100111;
		16'b0010111100111010: color_data = 12'b001110100111;
		16'b0010111100111011: color_data = 12'b001110100111;
		16'b0010111100111100: color_data = 12'b001110100111;
		16'b0010111100111101: color_data = 12'b001110100111;
		16'b0010111100111110: color_data = 12'b001110100111;
		16'b0010111100111111: color_data = 12'b001110100111;
		16'b0010111101000000: color_data = 12'b001110100111;
		16'b0010111101000001: color_data = 12'b001110100111;
		16'b0010111101000010: color_data = 12'b001110100111;
		16'b0010111101000011: color_data = 12'b001110100111;
		16'b0010111101000100: color_data = 12'b001110100111;
		16'b0010111101000101: color_data = 12'b001110100111;
		16'b0010111101000110: color_data = 12'b001110100111;
		16'b0010111101000111: color_data = 12'b001110100111;
		16'b0010111101001000: color_data = 12'b001110100111;
		16'b0010111101001001: color_data = 12'b001110100111;
		16'b0010111101001010: color_data = 12'b001110100111;
		16'b0010111101011110: color_data = 12'b001110100111;
		16'b0010111101011111: color_data = 12'b001110100111;
		16'b0010111101100000: color_data = 12'b001110100111;
		16'b0010111101100001: color_data = 12'b001110100111;
		16'b0010111101100010: color_data = 12'b001110100111;
		16'b0010111101100011: color_data = 12'b001110100111;
		16'b0010111101100100: color_data = 12'b001110100111;
		16'b0010111101100101: color_data = 12'b001110100111;
		16'b0010111101100110: color_data = 12'b001110100111;
		16'b0010111101100111: color_data = 12'b001110100111;
		16'b0010111101101000: color_data = 12'b001110100111;
		16'b0010111101101001: color_data = 12'b001110100111;
		16'b0010111101101010: color_data = 12'b001110100111;
		16'b0010111101101011: color_data = 12'b001110100111;
		16'b0010111101101100: color_data = 12'b001110100111;
		16'b0010111101101101: color_data = 12'b001110100111;
		16'b0010111101101110: color_data = 12'b001110100111;
		16'b0010111101101111: color_data = 12'b001110100111;
		16'b0010111101110000: color_data = 12'b001110100111;
		16'b0010111101110001: color_data = 12'b001110100111;
		16'b0010111101110010: color_data = 12'b001110100111;
		16'b0010111101110011: color_data = 12'b001110100111;
		16'b0010111101110100: color_data = 12'b001110100111;
		16'b0010111101110101: color_data = 12'b001110100111;
		16'b0010111101110110: color_data = 12'b001110100111;
		16'b0010111101110111: color_data = 12'b001110100111;
		16'b0010111101111000: color_data = 12'b001110100111;
		16'b0010111101111001: color_data = 12'b001110100111;
		16'b0010111101111010: color_data = 12'b001110100111;
		16'b0010111101111011: color_data = 12'b001110100111;
		16'b0011000000000111: color_data = 12'b001110100111;
		16'b0011000000001000: color_data = 12'b001110100111;
		16'b0011000000001001: color_data = 12'b001110100111;
		16'b0011000000001010: color_data = 12'b001110100111;
		16'b0011000000001011: color_data = 12'b001110100111;
		16'b0011000000001100: color_data = 12'b001110100111;
		16'b0011000000001101: color_data = 12'b001110100111;
		16'b0011000000001110: color_data = 12'b001110100111;
		16'b0011000000001111: color_data = 12'b001110100111;
		16'b0011000000010000: color_data = 12'b001110100111;
		16'b0011000000010001: color_data = 12'b001110100111;
		16'b0011000000010010: color_data = 12'b001110100111;
		16'b0011000000010011: color_data = 12'b001110100111;
		16'b0011000000010100: color_data = 12'b001110100111;
		16'b0011000000010101: color_data = 12'b001110100111;
		16'b0011000000010110: color_data = 12'b001110100111;
		16'b0011000000010111: color_data = 12'b001110100111;
		16'b0011000000011000: color_data = 12'b001110100111;
		16'b0011000000011001: color_data = 12'b001110100111;
		16'b0011000000011010: color_data = 12'b001110100111;
		16'b0011000000011011: color_data = 12'b001110100111;
		16'b0011000000011100: color_data = 12'b001110100111;
		16'b0011000000011101: color_data = 12'b001110100111;
		16'b0011000000011110: color_data = 12'b001110100111;
		16'b0011000000011111: color_data = 12'b001110100111;
		16'b0011000000100000: color_data = 12'b001110100111;
		16'b0011000000100001: color_data = 12'b001110100111;
		16'b0011000000100010: color_data = 12'b001110100111;
		16'b0011000000100011: color_data = 12'b001110100111;
		16'b0011000000100100: color_data = 12'b001110100111;
		16'b0011000000101011: color_data = 12'b001110100111;
		16'b0011000000101100: color_data = 12'b001110100111;
		16'b0011000000101101: color_data = 12'b001110100111;
		16'b0011000000101110: color_data = 12'b001110100111;
		16'b0011000000101111: color_data = 12'b001110100111;
		16'b0011000000110000: color_data = 12'b001110100111;
		16'b0011000000110001: color_data = 12'b001110100111;
		16'b0011000000110010: color_data = 12'b001110100111;
		16'b0011000000110011: color_data = 12'b001110100111;
		16'b0011000000110100: color_data = 12'b001110100111;
		16'b0011000000110101: color_data = 12'b001110100111;
		16'b0011000000110110: color_data = 12'b001110100111;
		16'b0011000000110111: color_data = 12'b001110100111;
		16'b0011000001000100: color_data = 12'b001110100111;
		16'b0011000001000101: color_data = 12'b001110100111;
		16'b0011000001000110: color_data = 12'b001110100111;
		16'b0011000001000111: color_data = 12'b001110100111;
		16'b0011000001001000: color_data = 12'b001110100111;
		16'b0011000001001001: color_data = 12'b001110100111;
		16'b0011000001001010: color_data = 12'b001110100111;
		16'b0011000001001011: color_data = 12'b001110100111;
		16'b0011000001001100: color_data = 12'b001110100111;
		16'b0011000001001101: color_data = 12'b001110100111;
		16'b0011000001001110: color_data = 12'b001110100111;
		16'b0011000001001111: color_data = 12'b001110100111;
		16'b0011000001010110: color_data = 12'b001110100111;
		16'b0011000001010111: color_data = 12'b001110100111;
		16'b0011000001011000: color_data = 12'b001110100111;
		16'b0011000001011001: color_data = 12'b001110100111;
		16'b0011000001011010: color_data = 12'b001110100111;
		16'b0011000001011011: color_data = 12'b001110100111;
		16'b0011000001011100: color_data = 12'b001110100111;
		16'b0011000001011101: color_data = 12'b001110100111;
		16'b0011000001011110: color_data = 12'b001110100111;
		16'b0011000001011111: color_data = 12'b001110100111;
		16'b0011000001100000: color_data = 12'b001110100111;
		16'b0011000001100001: color_data = 12'b001110100111;
		16'b0011000001100010: color_data = 12'b001110100111;
		16'b0011000001100011: color_data = 12'b001110100111;
		16'b0011000001100100: color_data = 12'b001110100111;
		16'b0011000001100101: color_data = 12'b001110100111;
		16'b0011000001100110: color_data = 12'b001110100111;
		16'b0011000001100111: color_data = 12'b001110100111;
		16'b0011000001101000: color_data = 12'b001110100111;
		16'b0011000001101001: color_data = 12'b001110100111;
		16'b0011000001101010: color_data = 12'b001110100111;
		16'b0011000001101011: color_data = 12'b001110100111;
		16'b0011000001101100: color_data = 12'b001110100111;
		16'b0011000001101101: color_data = 12'b001110100111;
		16'b0011000001101110: color_data = 12'b001110100111;
		16'b0011000001110101: color_data = 12'b001110100111;
		16'b0011000001110110: color_data = 12'b001110100111;
		16'b0011000001110111: color_data = 12'b001110100111;
		16'b0011000001111000: color_data = 12'b001110100111;
		16'b0011000001111001: color_data = 12'b001110100111;
		16'b0011000001111010: color_data = 12'b001110100111;
		16'b0011000001111011: color_data = 12'b001110100111;
		16'b0011000001111100: color_data = 12'b001110100111;
		16'b0011000001111101: color_data = 12'b001110100111;
		16'b0011000001111110: color_data = 12'b001110100111;
		16'b0011000001111111: color_data = 12'b001110100111;
		16'b0011000010000000: color_data = 12'b001110100111;
		16'b0011000010000001: color_data = 12'b001110100111;
		16'b0011000010000010: color_data = 12'b001110100111;
		16'b0011000010000011: color_data = 12'b001110100111;
		16'b0011000010000100: color_data = 12'b001110100111;
		16'b0011000010000101: color_data = 12'b001110100111;
		16'b0011000010000110: color_data = 12'b001110100111;
		16'b0011000010000111: color_data = 12'b001110100111;
		16'b0011000010001000: color_data = 12'b001110100111;
		16'b0011000010001001: color_data = 12'b001110100111;
		16'b0011000010001010: color_data = 12'b001110100111;
		16'b0011000010001011: color_data = 12'b001110100111;
		16'b0011000010001100: color_data = 12'b001110100111;
		16'b0011000010001101: color_data = 12'b001110100111;
		16'b0011000010001110: color_data = 12'b001110100111;
		16'b0011000010001111: color_data = 12'b001110100111;
		16'b0011000010010000: color_data = 12'b001110100111;
		16'b0011000010010001: color_data = 12'b001110100111;
		16'b0011000010010010: color_data = 12'b001110100111;
		16'b0011000010010011: color_data = 12'b001110100111;
		16'b0011000010100110: color_data = 12'b001110100111;
		16'b0011000010100111: color_data = 12'b001110100111;
		16'b0011000010101000: color_data = 12'b001110100111;
		16'b0011000010101001: color_data = 12'b001110100111;
		16'b0011000010101010: color_data = 12'b001110100111;
		16'b0011000010101011: color_data = 12'b001110100111;
		16'b0011000010101100: color_data = 12'b001110100111;
		16'b0011000010101101: color_data = 12'b001110100111;
		16'b0011000010101110: color_data = 12'b001110100111;
		16'b0011000010101111: color_data = 12'b001110100111;
		16'b0011000010110000: color_data = 12'b001110100111;
		16'b0011000010110001: color_data = 12'b001110100111;
		16'b0011000010110010: color_data = 12'b001110100111;
		16'b0011000010110011: color_data = 12'b001110100111;
		16'b0011000010110100: color_data = 12'b001110100111;
		16'b0011000010110101: color_data = 12'b001110100111;
		16'b0011000010110110: color_data = 12'b001110100111;
		16'b0011000010110111: color_data = 12'b001110100111;
		16'b0011000010111000: color_data = 12'b001110100111;
		16'b0011000010111001: color_data = 12'b001110100111;
		16'b0011000010111010: color_data = 12'b001110100111;
		16'b0011000010111011: color_data = 12'b001110100111;
		16'b0011000010111100: color_data = 12'b001110100111;
		16'b0011000010111101: color_data = 12'b001110100111;
		16'b0011000010111110: color_data = 12'b001110100111;
		16'b0011000010111111: color_data = 12'b001110100111;
		16'b0011000011000000: color_data = 12'b001110100111;
		16'b0011000011000001: color_data = 12'b001110100111;
		16'b0011000011000010: color_data = 12'b001110100111;
		16'b0011000011000011: color_data = 12'b001110100111;
		16'b0011000011000100: color_data = 12'b001110100111;
		16'b0011000011001011: color_data = 12'b001110100111;
		16'b0011000011001100: color_data = 12'b001110100111;
		16'b0011000011001101: color_data = 12'b001110100111;
		16'b0011000011001110: color_data = 12'b001110100111;
		16'b0011000011001111: color_data = 12'b001110100111;
		16'b0011000011010000: color_data = 12'b001110100111;
		16'b0011000011010001: color_data = 12'b001110100111;
		16'b0011000011010010: color_data = 12'b001110100111;
		16'b0011000011010011: color_data = 12'b001110100111;
		16'b0011000011010100: color_data = 12'b001110100111;
		16'b0011000011010101: color_data = 12'b001110100111;
		16'b0011000011010110: color_data = 12'b001110100111;
		16'b0011000011010111: color_data = 12'b001110100111;
		16'b0011000011011000: color_data = 12'b001110100111;
		16'b0011000011011001: color_data = 12'b001110100111;
		16'b0011000011011010: color_data = 12'b001110100111;
		16'b0011000011011011: color_data = 12'b001110100111;
		16'b0011000011011100: color_data = 12'b001110100111;
		16'b0011000011011101: color_data = 12'b001110100111;
		16'b0011000011011110: color_data = 12'b001110100111;
		16'b0011000011011111: color_data = 12'b001110100111;
		16'b0011000011100000: color_data = 12'b001110100111;
		16'b0011000011100001: color_data = 12'b001110100111;
		16'b0011000011100010: color_data = 12'b001110100111;
		16'b0011000011100011: color_data = 12'b001110100111;
		16'b0011000011100100: color_data = 12'b001110100111;
		16'b0011000011100101: color_data = 12'b001110100111;
		16'b0011000011100110: color_data = 12'b001110100111;
		16'b0011000011100111: color_data = 12'b001110100111;
		16'b0011000011101000: color_data = 12'b001110100111;
		16'b0011000011101001: color_data = 12'b001110100111;
		16'b0011000011101010: color_data = 12'b001110100111;
		16'b0011000011101011: color_data = 12'b001110100111;
		16'b0011000011101100: color_data = 12'b001110100111;
		16'b0011000011101101: color_data = 12'b001110100111;
		16'b0011000011101110: color_data = 12'b001110100111;
		16'b0011000011101111: color_data = 12'b001110100111;
		16'b0011000011110110: color_data = 12'b001110100111;
		16'b0011000011110111: color_data = 12'b001110100111;
		16'b0011000011111000: color_data = 12'b001110100111;
		16'b0011000011111001: color_data = 12'b001110100111;
		16'b0011000011111010: color_data = 12'b001110100111;
		16'b0011000011111011: color_data = 12'b001110100111;
		16'b0011000011111100: color_data = 12'b001110100111;
		16'b0011000011111101: color_data = 12'b001110100111;
		16'b0011000011111110: color_data = 12'b001110100111;
		16'b0011000011111111: color_data = 12'b001110100111;
		16'b0011000100000000: color_data = 12'b001110100111;
		16'b0011000100000001: color_data = 12'b001110100111;
		16'b0011000100000010: color_data = 12'b001110100111;
		16'b0011000100000011: color_data = 12'b001110100111;
		16'b0011000100000100: color_data = 12'b001110100111;
		16'b0011000100000101: color_data = 12'b001110100111;
		16'b0011000100000110: color_data = 12'b001110100111;
		16'b0011000100000111: color_data = 12'b001110100111;
		16'b0011000100001000: color_data = 12'b001110100111;
		16'b0011000100001001: color_data = 12'b001110100111;
		16'b0011000100001010: color_data = 12'b001110100111;
		16'b0011000100001011: color_data = 12'b001110100111;
		16'b0011000100001100: color_data = 12'b001110100111;
		16'b0011000100001101: color_data = 12'b001110100111;
		16'b0011000100001110: color_data = 12'b001110100111;
		16'b0011000100001111: color_data = 12'b001110100111;
		16'b0011000100010000: color_data = 12'b001110100111;
		16'b0011000100010001: color_data = 12'b001110100111;
		16'b0011000100010010: color_data = 12'b001110100111;
		16'b0011000100010011: color_data = 12'b001110100111;
		16'b0011000100010100: color_data = 12'b001110100111;
		16'b0011000100010101: color_data = 12'b001110100111;
		16'b0011000100010110: color_data = 12'b001110100111;
		16'b0011000100010111: color_data = 12'b001110100111;
		16'b0011000100011000: color_data = 12'b001110100111;
		16'b0011000100011001: color_data = 12'b001110100111;
		16'b0011000100011010: color_data = 12'b001110100111;
		16'b0011000100011011: color_data = 12'b001110100111;
		16'b0011000100011100: color_data = 12'b001110100111;
		16'b0011000100011101: color_data = 12'b001110100111;
		16'b0011000100011110: color_data = 12'b001110100111;
		16'b0011000100011111: color_data = 12'b001110100111;
		16'b0011000100100000: color_data = 12'b001110100111;
		16'b0011000100100001: color_data = 12'b001110100111;
		16'b0011000100100010: color_data = 12'b001110100111;
		16'b0011000100100011: color_data = 12'b001110100111;
		16'b0011000100100100: color_data = 12'b001110100111;
		16'b0011000100100101: color_data = 12'b001110100111;
		16'b0011000100100110: color_data = 12'b001110100111;
		16'b0011000100101101: color_data = 12'b001110100111;
		16'b0011000100101110: color_data = 12'b001110100111;
		16'b0011000100101111: color_data = 12'b001110100111;
		16'b0011000100110000: color_data = 12'b001110100111;
		16'b0011000100110001: color_data = 12'b001110100111;
		16'b0011000100110010: color_data = 12'b001110100111;
		16'b0011000100110011: color_data = 12'b001110100111;
		16'b0011000100110100: color_data = 12'b001110100111;
		16'b0011000100110101: color_data = 12'b001110100111;
		16'b0011000100110110: color_data = 12'b001110100111;
		16'b0011000100110111: color_data = 12'b001110100111;
		16'b0011000100111000: color_data = 12'b001110100111;
		16'b0011000100111001: color_data = 12'b001110100111;
		16'b0011000100111010: color_data = 12'b001110100111;
		16'b0011000100111011: color_data = 12'b001110100111;
		16'b0011000100111100: color_data = 12'b001110100111;
		16'b0011000100111101: color_data = 12'b001110100111;
		16'b0011000100111110: color_data = 12'b001110100111;
		16'b0011000100111111: color_data = 12'b001110100111;
		16'b0011000101000000: color_data = 12'b001110100111;
		16'b0011000101000001: color_data = 12'b001110100111;
		16'b0011000101000010: color_data = 12'b001110100111;
		16'b0011000101000011: color_data = 12'b001110100111;
		16'b0011000101000100: color_data = 12'b001110100111;
		16'b0011000101000101: color_data = 12'b001110100111;
		16'b0011000101000110: color_data = 12'b001110100111;
		16'b0011000101000111: color_data = 12'b001110100111;
		16'b0011000101001000: color_data = 12'b001110100111;
		16'b0011000101001001: color_data = 12'b001110100111;
		16'b0011000101001010: color_data = 12'b001110100111;
		16'b0011000101011110: color_data = 12'b001110100111;
		16'b0011000101011111: color_data = 12'b001110100111;
		16'b0011000101100000: color_data = 12'b001110100111;
		16'b0011000101100001: color_data = 12'b001110100111;
		16'b0011000101100010: color_data = 12'b001110100111;
		16'b0011000101100011: color_data = 12'b001110100111;
		16'b0011000101100100: color_data = 12'b001110100111;
		16'b0011000101100101: color_data = 12'b001110100111;
		16'b0011000101100110: color_data = 12'b001110100111;
		16'b0011000101100111: color_data = 12'b001110100111;
		16'b0011000101101000: color_data = 12'b001110100111;
		16'b0011000101101001: color_data = 12'b001110100111;
		16'b0011000101101010: color_data = 12'b001110100111;
		16'b0011000101101011: color_data = 12'b001110100111;
		16'b0011000101101100: color_data = 12'b001110100111;
		16'b0011000101101101: color_data = 12'b001110100111;
		16'b0011000101101110: color_data = 12'b001110100111;
		16'b0011000101101111: color_data = 12'b001110100111;
		16'b0011000101110000: color_data = 12'b001110100111;
		16'b0011000101110001: color_data = 12'b001110100111;
		16'b0011000101110010: color_data = 12'b001110100111;
		16'b0011000101110011: color_data = 12'b001110100111;
		16'b0011000101110100: color_data = 12'b001110100111;
		16'b0011000101110101: color_data = 12'b001110100111;
		16'b0011000101110110: color_data = 12'b001110100111;
		16'b0011000101110111: color_data = 12'b001110100111;
		16'b0011000101111000: color_data = 12'b001110100111;
		16'b0011000101111001: color_data = 12'b001110100111;
		16'b0011000101111010: color_data = 12'b001110100111;
		16'b0011000101111011: color_data = 12'b001110100111;
		16'b0011001000000111: color_data = 12'b001110100111;
		16'b0011001000001000: color_data = 12'b001110100111;
		16'b0011001000001001: color_data = 12'b001110100111;
		16'b0011001000001010: color_data = 12'b001110100111;
		16'b0011001000001011: color_data = 12'b001110100111;
		16'b0011001000001100: color_data = 12'b001110100111;
		16'b0011001000001101: color_data = 12'b001110100111;
		16'b0011001000001110: color_data = 12'b001110100111;
		16'b0011001000001111: color_data = 12'b001110100111;
		16'b0011001000010000: color_data = 12'b001110100111;
		16'b0011001000010001: color_data = 12'b001110100111;
		16'b0011001000010010: color_data = 12'b001110100111;
		16'b0011001000010011: color_data = 12'b001110100111;
		16'b0011001000010100: color_data = 12'b001110100111;
		16'b0011001000010101: color_data = 12'b001110100111;
		16'b0011001000010110: color_data = 12'b001110100111;
		16'b0011001000010111: color_data = 12'b001110100111;
		16'b0011001000011000: color_data = 12'b001110100111;
		16'b0011001000011001: color_data = 12'b001110100111;
		16'b0011001000011010: color_data = 12'b001110100111;
		16'b0011001000011011: color_data = 12'b001110100111;
		16'b0011001000011100: color_data = 12'b001110100111;
		16'b0011001000011101: color_data = 12'b001110100111;
		16'b0011001000011110: color_data = 12'b001110100111;
		16'b0011001000011111: color_data = 12'b001110100111;
		16'b0011001000100000: color_data = 12'b001110100111;
		16'b0011001000100001: color_data = 12'b001110100111;
		16'b0011001000100010: color_data = 12'b001110100111;
		16'b0011001000100011: color_data = 12'b001110100111;
		16'b0011001000100100: color_data = 12'b001110100111;
		16'b0011001000101011: color_data = 12'b001110100111;
		16'b0011001000101100: color_data = 12'b001110100111;
		16'b0011001000101101: color_data = 12'b001110100111;
		16'b0011001000101110: color_data = 12'b001110100111;
		16'b0011001000101111: color_data = 12'b001110100111;
		16'b0011001000110000: color_data = 12'b001110100111;
		16'b0011001000110001: color_data = 12'b001110100111;
		16'b0011001000110010: color_data = 12'b001110100111;
		16'b0011001000110011: color_data = 12'b001110100111;
		16'b0011001000110100: color_data = 12'b001110100111;
		16'b0011001000110101: color_data = 12'b001110100111;
		16'b0011001000110110: color_data = 12'b001110100111;
		16'b0011001000110111: color_data = 12'b001110100111;
		16'b0011001001000100: color_data = 12'b001110100111;
		16'b0011001001000101: color_data = 12'b001110100111;
		16'b0011001001000110: color_data = 12'b001110100111;
		16'b0011001001000111: color_data = 12'b001110100111;
		16'b0011001001001000: color_data = 12'b001110100111;
		16'b0011001001001001: color_data = 12'b001110100111;
		16'b0011001001001010: color_data = 12'b001110100111;
		16'b0011001001001011: color_data = 12'b001110100111;
		16'b0011001001001100: color_data = 12'b001110100111;
		16'b0011001001001101: color_data = 12'b001110100111;
		16'b0011001001001110: color_data = 12'b001110100111;
		16'b0011001001001111: color_data = 12'b001110100111;
		16'b0011001001010110: color_data = 12'b001110100111;
		16'b0011001001010111: color_data = 12'b001110100111;
		16'b0011001001011000: color_data = 12'b001110100111;
		16'b0011001001011001: color_data = 12'b001110100111;
		16'b0011001001011010: color_data = 12'b001110100111;
		16'b0011001001011011: color_data = 12'b001110100111;
		16'b0011001001011100: color_data = 12'b001110100111;
		16'b0011001001011101: color_data = 12'b001110100111;
		16'b0011001001011110: color_data = 12'b001110100111;
		16'b0011001001011111: color_data = 12'b001110100111;
		16'b0011001001100000: color_data = 12'b001110100111;
		16'b0011001001100001: color_data = 12'b001110100111;
		16'b0011001001100010: color_data = 12'b001110100111;
		16'b0011001001100011: color_data = 12'b001110100111;
		16'b0011001001100100: color_data = 12'b001110100111;
		16'b0011001001100101: color_data = 12'b001110100111;
		16'b0011001001100110: color_data = 12'b001110100111;
		16'b0011001001100111: color_data = 12'b001110100111;
		16'b0011001001101000: color_data = 12'b001110100111;
		16'b0011001001101001: color_data = 12'b001110100111;
		16'b0011001001101010: color_data = 12'b001110100111;
		16'b0011001001101011: color_data = 12'b001110100111;
		16'b0011001001101100: color_data = 12'b001110100111;
		16'b0011001001101101: color_data = 12'b001110100111;
		16'b0011001001101110: color_data = 12'b001110100111;
		16'b0011001001110101: color_data = 12'b001110100111;
		16'b0011001001110110: color_data = 12'b001110100111;
		16'b0011001001110111: color_data = 12'b001110100111;
		16'b0011001001111000: color_data = 12'b001110100111;
		16'b0011001001111001: color_data = 12'b001110100111;
		16'b0011001001111010: color_data = 12'b001110100111;
		16'b0011001001111011: color_data = 12'b001110100111;
		16'b0011001001111100: color_data = 12'b001110100111;
		16'b0011001001111101: color_data = 12'b001110100111;
		16'b0011001001111110: color_data = 12'b001110100111;
		16'b0011001001111111: color_data = 12'b001110100111;
		16'b0011001010000000: color_data = 12'b001110100111;
		16'b0011001010000001: color_data = 12'b001110100111;
		16'b0011001010000010: color_data = 12'b001110100111;
		16'b0011001010000011: color_data = 12'b001110100111;
		16'b0011001010000100: color_data = 12'b001110100111;
		16'b0011001010000101: color_data = 12'b001110100111;
		16'b0011001010000110: color_data = 12'b001110100111;
		16'b0011001010000111: color_data = 12'b001110100111;
		16'b0011001010001000: color_data = 12'b001110100111;
		16'b0011001010001001: color_data = 12'b001110100111;
		16'b0011001010001010: color_data = 12'b001110100111;
		16'b0011001010001011: color_data = 12'b001110100111;
		16'b0011001010001100: color_data = 12'b001110100111;
		16'b0011001010001101: color_data = 12'b001110100111;
		16'b0011001010001110: color_data = 12'b001110100111;
		16'b0011001010001111: color_data = 12'b001110100111;
		16'b0011001010010000: color_data = 12'b001110100111;
		16'b0011001010010001: color_data = 12'b001110100111;
		16'b0011001010010010: color_data = 12'b001110100111;
		16'b0011001010010011: color_data = 12'b001110100111;
		16'b0011001010100110: color_data = 12'b001110100111;
		16'b0011001010100111: color_data = 12'b001110100111;
		16'b0011001010101000: color_data = 12'b001110100111;
		16'b0011001010101001: color_data = 12'b001110100111;
		16'b0011001010101010: color_data = 12'b001110100111;
		16'b0011001010101011: color_data = 12'b001110100111;
		16'b0011001010101100: color_data = 12'b001110100111;
		16'b0011001010101101: color_data = 12'b001110100111;
		16'b0011001010101110: color_data = 12'b001110100111;
		16'b0011001010101111: color_data = 12'b001110100111;
		16'b0011001010110000: color_data = 12'b001110100111;
		16'b0011001010110001: color_data = 12'b001110100111;
		16'b0011001010110010: color_data = 12'b001110100111;
		16'b0011001010110011: color_data = 12'b001110100111;
		16'b0011001010110100: color_data = 12'b001110100111;
		16'b0011001010110101: color_data = 12'b001110100111;
		16'b0011001010110110: color_data = 12'b001110100111;
		16'b0011001010110111: color_data = 12'b001110100111;
		16'b0011001010111000: color_data = 12'b001110100111;
		16'b0011001010111001: color_data = 12'b001110100111;
		16'b0011001010111010: color_data = 12'b001110100111;
		16'b0011001010111011: color_data = 12'b001110100111;
		16'b0011001010111100: color_data = 12'b001110100111;
		16'b0011001010111101: color_data = 12'b001110100111;
		16'b0011001010111110: color_data = 12'b001110100111;
		16'b0011001010111111: color_data = 12'b001110100111;
		16'b0011001011000000: color_data = 12'b001110100111;
		16'b0011001011000001: color_data = 12'b001110100111;
		16'b0011001011000010: color_data = 12'b001110100111;
		16'b0011001011000011: color_data = 12'b001110100111;
		16'b0011001011000100: color_data = 12'b001110100111;
		16'b0011001011001011: color_data = 12'b001110100111;
		16'b0011001011001100: color_data = 12'b001110100111;
		16'b0011001011001101: color_data = 12'b001110100111;
		16'b0011001011001110: color_data = 12'b001110100111;
		16'b0011001011001111: color_data = 12'b001110100111;
		16'b0011001011010000: color_data = 12'b001110100111;
		16'b0011001011010001: color_data = 12'b001110100111;
		16'b0011001011010010: color_data = 12'b001110100111;
		16'b0011001011010011: color_data = 12'b001110100111;
		16'b0011001011010100: color_data = 12'b001110100111;
		16'b0011001011010101: color_data = 12'b001110100111;
		16'b0011001011010110: color_data = 12'b001110100111;
		16'b0011001011010111: color_data = 12'b001110100111;
		16'b0011001011011000: color_data = 12'b001110100111;
		16'b0011001011011001: color_data = 12'b001110100111;
		16'b0011001011011010: color_data = 12'b001110100111;
		16'b0011001011011011: color_data = 12'b001110100111;
		16'b0011001011011100: color_data = 12'b001110100111;
		16'b0011001011011101: color_data = 12'b001110100111;
		16'b0011001011011110: color_data = 12'b001110100111;
		16'b0011001011011111: color_data = 12'b001110100111;
		16'b0011001011100000: color_data = 12'b001110100111;
		16'b0011001011100001: color_data = 12'b001110100111;
		16'b0011001011100010: color_data = 12'b001110100111;
		16'b0011001011100011: color_data = 12'b001110100111;
		16'b0011001011100100: color_data = 12'b001110100111;
		16'b0011001011100101: color_data = 12'b001110100111;
		16'b0011001011100110: color_data = 12'b001110100111;
		16'b0011001011100111: color_data = 12'b001110100111;
		16'b0011001011101000: color_data = 12'b001110100111;
		16'b0011001011101001: color_data = 12'b001110100111;
		16'b0011001011101010: color_data = 12'b001110100111;
		16'b0011001011101011: color_data = 12'b001110100111;
		16'b0011001011101100: color_data = 12'b001110100111;
		16'b0011001011101101: color_data = 12'b001110100111;
		16'b0011001011101110: color_data = 12'b001110100111;
		16'b0011001011101111: color_data = 12'b001110100111;
		16'b0011001011110110: color_data = 12'b001110100111;
		16'b0011001011110111: color_data = 12'b001110100111;
		16'b0011001011111000: color_data = 12'b001110100111;
		16'b0011001011111001: color_data = 12'b001110100111;
		16'b0011001011111010: color_data = 12'b001110100111;
		16'b0011001011111011: color_data = 12'b001110100111;
		16'b0011001011111100: color_data = 12'b001110100111;
		16'b0011001011111101: color_data = 12'b001110100111;
		16'b0011001011111110: color_data = 12'b001110100111;
		16'b0011001011111111: color_data = 12'b001110100111;
		16'b0011001100000000: color_data = 12'b001110100111;
		16'b0011001100000001: color_data = 12'b001110100111;
		16'b0011001100000010: color_data = 12'b001110100111;
		16'b0011001100000011: color_data = 12'b001110100111;
		16'b0011001100000100: color_data = 12'b001110100111;
		16'b0011001100000101: color_data = 12'b001110100111;
		16'b0011001100000110: color_data = 12'b001110100111;
		16'b0011001100000111: color_data = 12'b001110100111;
		16'b0011001100001000: color_data = 12'b001110100111;
		16'b0011001100001001: color_data = 12'b001110100111;
		16'b0011001100001010: color_data = 12'b001110100111;
		16'b0011001100001011: color_data = 12'b001110100111;
		16'b0011001100001100: color_data = 12'b001110100111;
		16'b0011001100001101: color_data = 12'b001110100111;
		16'b0011001100001110: color_data = 12'b001110100111;
		16'b0011001100001111: color_data = 12'b001110100111;
		16'b0011001100010000: color_data = 12'b001110100111;
		16'b0011001100010001: color_data = 12'b001110100111;
		16'b0011001100010010: color_data = 12'b001110100111;
		16'b0011001100010011: color_data = 12'b001110100111;
		16'b0011001100010100: color_data = 12'b001110100111;
		16'b0011001100010101: color_data = 12'b001110100111;
		16'b0011001100010110: color_data = 12'b001110100111;
		16'b0011001100010111: color_data = 12'b001110100111;
		16'b0011001100011000: color_data = 12'b001110100111;
		16'b0011001100011001: color_data = 12'b001110100111;
		16'b0011001100011010: color_data = 12'b001110100111;
		16'b0011001100011011: color_data = 12'b001110100111;
		16'b0011001100011100: color_data = 12'b001110100111;
		16'b0011001100011101: color_data = 12'b001110100111;
		16'b0011001100011110: color_data = 12'b001110100111;
		16'b0011001100011111: color_data = 12'b001110100111;
		16'b0011001100100000: color_data = 12'b001110100111;
		16'b0011001100100001: color_data = 12'b001110100111;
		16'b0011001100100010: color_data = 12'b001110100111;
		16'b0011001100100011: color_data = 12'b001110100111;
		16'b0011001100100100: color_data = 12'b001110100111;
		16'b0011001100100101: color_data = 12'b001110100111;
		16'b0011001100100110: color_data = 12'b001110100111;
		16'b0011001100101101: color_data = 12'b001110100111;
		16'b0011001100101110: color_data = 12'b001110100111;
		16'b0011001100101111: color_data = 12'b001110100111;
		16'b0011001100110000: color_data = 12'b001110100111;
		16'b0011001100110001: color_data = 12'b001110100111;
		16'b0011001100110010: color_data = 12'b001110100111;
		16'b0011001100110011: color_data = 12'b001110100111;
		16'b0011001100110100: color_data = 12'b001110100111;
		16'b0011001100110101: color_data = 12'b001110100111;
		16'b0011001100110110: color_data = 12'b001110100111;
		16'b0011001100110111: color_data = 12'b001110100111;
		16'b0011001100111000: color_data = 12'b001110100111;
		16'b0011001100111001: color_data = 12'b001110100111;
		16'b0011001100111010: color_data = 12'b001110100111;
		16'b0011001100111011: color_data = 12'b001110100111;
		16'b0011001100111100: color_data = 12'b001110100111;
		16'b0011001100111101: color_data = 12'b001110100111;
		16'b0011001100111110: color_data = 12'b001110100111;
		16'b0011001100111111: color_data = 12'b001110100111;
		16'b0011001101000000: color_data = 12'b001110100111;
		16'b0011001101000001: color_data = 12'b001110100111;
		16'b0011001101000010: color_data = 12'b001110100111;
		16'b0011001101000011: color_data = 12'b001110100111;
		16'b0011001101000100: color_data = 12'b001110100111;
		16'b0011001101000101: color_data = 12'b001110100111;
		16'b0011001101000110: color_data = 12'b001110100111;
		16'b0011001101000111: color_data = 12'b001110100111;
		16'b0011001101001000: color_data = 12'b001110100111;
		16'b0011001101001001: color_data = 12'b001110100111;
		16'b0011001101001010: color_data = 12'b001110100111;
		16'b0011001101011110: color_data = 12'b001110100111;
		16'b0011001101011111: color_data = 12'b001110100111;
		16'b0011001101100000: color_data = 12'b001110100111;
		16'b0011001101100001: color_data = 12'b001110100111;
		16'b0011001101100010: color_data = 12'b001110100111;
		16'b0011001101100011: color_data = 12'b001110100111;
		16'b0011001101100100: color_data = 12'b001110100111;
		16'b0011001101100101: color_data = 12'b001110100111;
		16'b0011001101100110: color_data = 12'b001110100111;
		16'b0011001101100111: color_data = 12'b001110100111;
		16'b0011001101101000: color_data = 12'b001110100111;
		16'b0011001101101001: color_data = 12'b001110100111;
		16'b0011001101101010: color_data = 12'b001110100111;
		16'b0011001101101011: color_data = 12'b001110100111;
		16'b0011001101101100: color_data = 12'b001110100111;
		16'b0011001101101101: color_data = 12'b001110100111;
		16'b0011001101101110: color_data = 12'b001110100111;
		16'b0011001101101111: color_data = 12'b001110100111;
		16'b0011001101110000: color_data = 12'b001110100111;
		16'b0011001101110001: color_data = 12'b001110100111;
		16'b0011001101110010: color_data = 12'b001110100111;
		16'b0011001101110011: color_data = 12'b001110100111;
		16'b0011001101110100: color_data = 12'b001110100111;
		16'b0011001101110101: color_data = 12'b001110100111;
		16'b0011001101110110: color_data = 12'b001110100111;
		16'b0011001101110111: color_data = 12'b001110100111;
		16'b0011001101111000: color_data = 12'b001110100111;
		16'b0011001101111001: color_data = 12'b001110100111;
		16'b0011001101111010: color_data = 12'b001110100111;
		16'b0011001101111011: color_data = 12'b001110100111;
		16'b0011010000000000: color_data = 12'b001110100111;
		16'b0011010000000001: color_data = 12'b001110100111;
		16'b0011010000000010: color_data = 12'b001110100111;
		16'b0011010000000011: color_data = 12'b001110100111;
		16'b0011010000000100: color_data = 12'b001110100111;
		16'b0011010000000101: color_data = 12'b001110100111;
		16'b0011010000000110: color_data = 12'b001110100111;
		16'b0011010000000111: color_data = 12'b001110100111;
		16'b0011010000001000: color_data = 12'b001110100111;
		16'b0011010000001001: color_data = 12'b001110100111;
		16'b0011010000001010: color_data = 12'b001110100111;
		16'b0011010000001011: color_data = 12'b001110100111;
		16'b0011010000001100: color_data = 12'b001110100111;
		16'b0011010000001101: color_data = 12'b001110100111;
		16'b0011010000001110: color_data = 12'b001110100111;
		16'b0011010000001111: color_data = 12'b001110100111;
		16'b0011010000010000: color_data = 12'b001110100111;
		16'b0011010000010001: color_data = 12'b001110100111;
		16'b0011010000010010: color_data = 12'b001110100111;
		16'b0011010000101011: color_data = 12'b001110100111;
		16'b0011010000101100: color_data = 12'b001110100111;
		16'b0011010000101101: color_data = 12'b001110100111;
		16'b0011010000101110: color_data = 12'b001110100111;
		16'b0011010000101111: color_data = 12'b001110100111;
		16'b0011010000110000: color_data = 12'b001110100111;
		16'b0011010000110001: color_data = 12'b001110100111;
		16'b0011010000110010: color_data = 12'b001110100111;
		16'b0011010000110011: color_data = 12'b001110100111;
		16'b0011010000110100: color_data = 12'b001110100111;
		16'b0011010000110101: color_data = 12'b001110100111;
		16'b0011010000110110: color_data = 12'b001110100111;
		16'b0011010000110111: color_data = 12'b001110100111;
		16'b0011010001000100: color_data = 12'b001110100111;
		16'b0011010001000101: color_data = 12'b001110100111;
		16'b0011010001000110: color_data = 12'b001110100111;
		16'b0011010001000111: color_data = 12'b001110100111;
		16'b0011010001001000: color_data = 12'b001110100111;
		16'b0011010001001001: color_data = 12'b001110100111;
		16'b0011010001001010: color_data = 12'b001110100111;
		16'b0011010001001011: color_data = 12'b001110100111;
		16'b0011010001001100: color_data = 12'b001110100111;
		16'b0011010001001101: color_data = 12'b001110100111;
		16'b0011010001001110: color_data = 12'b001110100111;
		16'b0011010001001111: color_data = 12'b001110100111;
		16'b0011010001011100: color_data = 12'b001110100111;
		16'b0011010001011101: color_data = 12'b001110100111;
		16'b0011010001011110: color_data = 12'b001110100111;
		16'b0011010001011111: color_data = 12'b001110100111;
		16'b0011010001100000: color_data = 12'b001110100111;
		16'b0011010001100001: color_data = 12'b001110100111;
		16'b0011010001100010: color_data = 12'b001110100111;
		16'b0011010001100011: color_data = 12'b001110100111;
		16'b0011010001100100: color_data = 12'b001110100111;
		16'b0011010001100101: color_data = 12'b001110100111;
		16'b0011010001100110: color_data = 12'b001110100111;
		16'b0011010001100111: color_data = 12'b001110100111;
		16'b0011010001101000: color_data = 12'b001110100111;
		16'b0011010001110101: color_data = 12'b001110100111;
		16'b0011010001110110: color_data = 12'b001110100111;
		16'b0011010001110111: color_data = 12'b001110100111;
		16'b0011010001111000: color_data = 12'b001110100111;
		16'b0011010001111001: color_data = 12'b001110100111;
		16'b0011010001111010: color_data = 12'b001110100111;
		16'b0011010001111011: color_data = 12'b001110100111;
		16'b0011010001111100: color_data = 12'b001110100111;
		16'b0011010001111101: color_data = 12'b001110100111;
		16'b0011010001111110: color_data = 12'b001110100111;
		16'b0011010001111111: color_data = 12'b001110100111;
		16'b0011010010000000: color_data = 12'b001110100111;
		16'b0011010010001101: color_data = 12'b001110100111;
		16'b0011010010001110: color_data = 12'b001110100111;
		16'b0011010010001111: color_data = 12'b001110100111;
		16'b0011010010010000: color_data = 12'b001110100111;
		16'b0011010010010001: color_data = 12'b001110100111;
		16'b0011010010010010: color_data = 12'b001110100111;
		16'b0011010010010011: color_data = 12'b001110100111;
		16'b0011010010010100: color_data = 12'b001110100111;
		16'b0011010010010101: color_data = 12'b001110100111;
		16'b0011010010010110: color_data = 12'b001110100111;
		16'b0011010010010111: color_data = 12'b001110100111;
		16'b0011010010011000: color_data = 12'b001110100111;
		16'b0011010010011001: color_data = 12'b001110100111;
		16'b0011010010100000: color_data = 12'b001110100111;
		16'b0011010010100001: color_data = 12'b001110100111;
		16'b0011010010100010: color_data = 12'b001110100111;
		16'b0011010010100011: color_data = 12'b001110100111;
		16'b0011010010100100: color_data = 12'b001110100111;
		16'b0011010010100101: color_data = 12'b001110100111;
		16'b0011010010100110: color_data = 12'b001110100111;
		16'b0011010010100111: color_data = 12'b001110100111;
		16'b0011010010101000: color_data = 12'b001110100111;
		16'b0011010010101001: color_data = 12'b001110100111;
		16'b0011010010101010: color_data = 12'b001110100111;
		16'b0011010010101011: color_data = 12'b001110100111;
		16'b0011010011001011: color_data = 12'b001110100111;
		16'b0011010011001100: color_data = 12'b001110100111;
		16'b0011010011001101: color_data = 12'b001110100111;
		16'b0011010011001110: color_data = 12'b001110100111;
		16'b0011010011001111: color_data = 12'b001110100111;
		16'b0011010011010000: color_data = 12'b001110100111;
		16'b0011010011010001: color_data = 12'b001110100111;
		16'b0011010011010010: color_data = 12'b001110100111;
		16'b0011010011010011: color_data = 12'b001110100111;
		16'b0011010011010100: color_data = 12'b001110100111;
		16'b0011010011010101: color_data = 12'b001110100111;
		16'b0011010011010110: color_data = 12'b001110100111;
		16'b0011010011100011: color_data = 12'b001110100111;
		16'b0011010011100100: color_data = 12'b001110100111;
		16'b0011010011100101: color_data = 12'b001110100111;
		16'b0011010011100110: color_data = 12'b001110100111;
		16'b0011010011100111: color_data = 12'b001110100111;
		16'b0011010011101000: color_data = 12'b001110100111;
		16'b0011010011101001: color_data = 12'b001110100111;
		16'b0011010011101010: color_data = 12'b001110100111;
		16'b0011010011101011: color_data = 12'b001110100111;
		16'b0011010011101100: color_data = 12'b001110100111;
		16'b0011010011101101: color_data = 12'b001110100111;
		16'b0011010011101110: color_data = 12'b001110100111;
		16'b0011010011101111: color_data = 12'b001110100111;
		16'b0011010011110110: color_data = 12'b001110100111;
		16'b0011010011110111: color_data = 12'b001110100111;
		16'b0011010011111000: color_data = 12'b001110100111;
		16'b0011010011111001: color_data = 12'b001110100111;
		16'b0011010011111010: color_data = 12'b001110100111;
		16'b0011010011111011: color_data = 12'b001110100111;
		16'b0011010011111100: color_data = 12'b001110100111;
		16'b0011010011111101: color_data = 12'b001110100111;
		16'b0011010011111110: color_data = 12'b001110100111;
		16'b0011010011111111: color_data = 12'b001110100111;
		16'b0011010100000000: color_data = 12'b001110100111;
		16'b0011010100000001: color_data = 12'b001110100111;
		16'b0011010100011010: color_data = 12'b001110100111;
		16'b0011010100011011: color_data = 12'b001110100111;
		16'b0011010100011100: color_data = 12'b001110100111;
		16'b0011010100011101: color_data = 12'b001110100111;
		16'b0011010100011110: color_data = 12'b001110100111;
		16'b0011010100011111: color_data = 12'b001110100111;
		16'b0011010100100000: color_data = 12'b001110100111;
		16'b0011010100100001: color_data = 12'b001110100111;
		16'b0011010100100010: color_data = 12'b001110100111;
		16'b0011010100100011: color_data = 12'b001110100111;
		16'b0011010100100100: color_data = 12'b001110100111;
		16'b0011010100100101: color_data = 12'b001110100111;
		16'b0011010100100110: color_data = 12'b001110100111;
		16'b0011010100101101: color_data = 12'b001110100111;
		16'b0011010100101110: color_data = 12'b001110100111;
		16'b0011010100101111: color_data = 12'b001110100111;
		16'b0011010100110000: color_data = 12'b001110100111;
		16'b0011010100110001: color_data = 12'b001110100111;
		16'b0011010100110010: color_data = 12'b001110100111;
		16'b0011010100110011: color_data = 12'b001110100111;
		16'b0011010100110100: color_data = 12'b001110100111;
		16'b0011010100110101: color_data = 12'b001110100111;
		16'b0011010100110110: color_data = 12'b001110100111;
		16'b0011010100110111: color_data = 12'b001110100111;
		16'b0011010100111000: color_data = 12'b001110100111;
		16'b0011010101000101: color_data = 12'b001110100111;
		16'b0011010101000110: color_data = 12'b001110100111;
		16'b0011010101000111: color_data = 12'b001110100111;
		16'b0011010101001000: color_data = 12'b001110100111;
		16'b0011010101001001: color_data = 12'b001110100111;
		16'b0011010101001010: color_data = 12'b001110100111;
		16'b0011010101001011: color_data = 12'b001110100111;
		16'b0011010101001100: color_data = 12'b001110100111;
		16'b0011010101001101: color_data = 12'b001110100111;
		16'b0011010101001110: color_data = 12'b001110100111;
		16'b0011010101001111: color_data = 12'b001110100111;
		16'b0011010101010000: color_data = 12'b001110100111;
		16'b0011010101010001: color_data = 12'b001110100111;
		16'b0011010101011000: color_data = 12'b001110100111;
		16'b0011010101011001: color_data = 12'b001110100111;
		16'b0011010101011010: color_data = 12'b001110100111;
		16'b0011010101011011: color_data = 12'b001110100111;
		16'b0011010101011100: color_data = 12'b001110100111;
		16'b0011010101011101: color_data = 12'b001110100111;
		16'b0011010101011110: color_data = 12'b001110100111;
		16'b0011010101011111: color_data = 12'b001110100111;
		16'b0011010101100000: color_data = 12'b001110100111;
		16'b0011010101100001: color_data = 12'b001110100111;
		16'b0011010101100010: color_data = 12'b001110100111;
		16'b0011010101100011: color_data = 12'b001110100111;
		16'b0011011000000000: color_data = 12'b001110100111;
		16'b0011011000000001: color_data = 12'b001110100111;
		16'b0011011000000010: color_data = 12'b001110100111;
		16'b0011011000000011: color_data = 12'b001110100111;
		16'b0011011000000100: color_data = 12'b001110100111;
		16'b0011011000000101: color_data = 12'b001110100111;
		16'b0011011000000110: color_data = 12'b001110100111;
		16'b0011011000000111: color_data = 12'b001110100111;
		16'b0011011000001000: color_data = 12'b001110100111;
		16'b0011011000001001: color_data = 12'b001110100111;
		16'b0011011000001010: color_data = 12'b001110100111;
		16'b0011011000001011: color_data = 12'b001110100111;
		16'b0011011000001100: color_data = 12'b001110100111;
		16'b0011011000001101: color_data = 12'b001110100111;
		16'b0011011000001110: color_data = 12'b001110100111;
		16'b0011011000001111: color_data = 12'b001110100111;
		16'b0011011000010000: color_data = 12'b001110100111;
		16'b0011011000010001: color_data = 12'b001110100111;
		16'b0011011000010010: color_data = 12'b001110100111;
		16'b0011011000101011: color_data = 12'b001110100111;
		16'b0011011000101100: color_data = 12'b001110100111;
		16'b0011011000101101: color_data = 12'b001110100111;
		16'b0011011000101110: color_data = 12'b001110100111;
		16'b0011011000101111: color_data = 12'b001110100111;
		16'b0011011000110000: color_data = 12'b001110100111;
		16'b0011011000110001: color_data = 12'b001110100111;
		16'b0011011000110010: color_data = 12'b001110100111;
		16'b0011011000110011: color_data = 12'b001110100111;
		16'b0011011000110100: color_data = 12'b001110100111;
		16'b0011011000110101: color_data = 12'b001110100111;
		16'b0011011000110110: color_data = 12'b001110100111;
		16'b0011011000110111: color_data = 12'b001110100111;
		16'b0011011001000100: color_data = 12'b001110100111;
		16'b0011011001000101: color_data = 12'b001110100111;
		16'b0011011001000110: color_data = 12'b001110100111;
		16'b0011011001000111: color_data = 12'b001110100111;
		16'b0011011001001000: color_data = 12'b001110100111;
		16'b0011011001001001: color_data = 12'b001110100111;
		16'b0011011001001010: color_data = 12'b001110100111;
		16'b0011011001001011: color_data = 12'b001110100111;
		16'b0011011001001100: color_data = 12'b001110100111;
		16'b0011011001001101: color_data = 12'b001110100111;
		16'b0011011001001110: color_data = 12'b001110100111;
		16'b0011011001001111: color_data = 12'b001110100111;
		16'b0011011001011100: color_data = 12'b001110100111;
		16'b0011011001011101: color_data = 12'b001110100111;
		16'b0011011001011110: color_data = 12'b001110100111;
		16'b0011011001011111: color_data = 12'b001110100111;
		16'b0011011001100000: color_data = 12'b001110100111;
		16'b0011011001100001: color_data = 12'b001110100111;
		16'b0011011001100010: color_data = 12'b001110100111;
		16'b0011011001100011: color_data = 12'b001110100111;
		16'b0011011001100100: color_data = 12'b001110100111;
		16'b0011011001100101: color_data = 12'b001110100111;
		16'b0011011001100110: color_data = 12'b001110100111;
		16'b0011011001100111: color_data = 12'b001110100111;
		16'b0011011001101000: color_data = 12'b001110100111;
		16'b0011011001110101: color_data = 12'b001110100111;
		16'b0011011001110110: color_data = 12'b001110100111;
		16'b0011011001110111: color_data = 12'b001110100111;
		16'b0011011001111000: color_data = 12'b001110100111;
		16'b0011011001111001: color_data = 12'b001110100111;
		16'b0011011001111010: color_data = 12'b001110100111;
		16'b0011011001111011: color_data = 12'b001110100111;
		16'b0011011001111100: color_data = 12'b001110100111;
		16'b0011011001111101: color_data = 12'b001110100111;
		16'b0011011001111110: color_data = 12'b001110100111;
		16'b0011011001111111: color_data = 12'b001110100111;
		16'b0011011010000000: color_data = 12'b001110100111;
		16'b0011011010001101: color_data = 12'b001110100111;
		16'b0011011010001110: color_data = 12'b001110100111;
		16'b0011011010001111: color_data = 12'b001110100111;
		16'b0011011010010000: color_data = 12'b001110100111;
		16'b0011011010010001: color_data = 12'b001110100111;
		16'b0011011010010010: color_data = 12'b001110100111;
		16'b0011011010010011: color_data = 12'b001110100111;
		16'b0011011010010100: color_data = 12'b001110100111;
		16'b0011011010010101: color_data = 12'b001110100111;
		16'b0011011010010110: color_data = 12'b001110100111;
		16'b0011011010010111: color_data = 12'b001110100111;
		16'b0011011010011000: color_data = 12'b001110100111;
		16'b0011011010011001: color_data = 12'b001110100111;
		16'b0011011010100000: color_data = 12'b001110100111;
		16'b0011011010100001: color_data = 12'b001110100111;
		16'b0011011010100010: color_data = 12'b001110100111;
		16'b0011011010100011: color_data = 12'b001110100111;
		16'b0011011010100100: color_data = 12'b001110100111;
		16'b0011011010100101: color_data = 12'b001110100111;
		16'b0011011010100110: color_data = 12'b001110100111;
		16'b0011011010100111: color_data = 12'b001110100111;
		16'b0011011010101000: color_data = 12'b001110100111;
		16'b0011011010101001: color_data = 12'b001110100111;
		16'b0011011010101010: color_data = 12'b001110100111;
		16'b0011011010101011: color_data = 12'b001110100111;
		16'b0011011011001011: color_data = 12'b001110100111;
		16'b0011011011001100: color_data = 12'b001110100111;
		16'b0011011011001101: color_data = 12'b001110100111;
		16'b0011011011001110: color_data = 12'b001110100111;
		16'b0011011011001111: color_data = 12'b001110100111;
		16'b0011011011010000: color_data = 12'b001110100111;
		16'b0011011011010001: color_data = 12'b001110100111;
		16'b0011011011010010: color_data = 12'b001110100111;
		16'b0011011011010011: color_data = 12'b001110100111;
		16'b0011011011010100: color_data = 12'b001110100111;
		16'b0011011011010101: color_data = 12'b001110100111;
		16'b0011011011010110: color_data = 12'b001110100111;
		16'b0011011011100011: color_data = 12'b001110100111;
		16'b0011011011100100: color_data = 12'b001110100111;
		16'b0011011011100101: color_data = 12'b001110100111;
		16'b0011011011100110: color_data = 12'b001110100111;
		16'b0011011011100111: color_data = 12'b001110100111;
		16'b0011011011101000: color_data = 12'b001110100111;
		16'b0011011011101001: color_data = 12'b001110100111;
		16'b0011011011101010: color_data = 12'b001110100111;
		16'b0011011011101011: color_data = 12'b001110100111;
		16'b0011011011101100: color_data = 12'b001110100111;
		16'b0011011011101101: color_data = 12'b001110100111;
		16'b0011011011101110: color_data = 12'b001110100111;
		16'b0011011011101111: color_data = 12'b001110100111;
		16'b0011011011110110: color_data = 12'b001110100111;
		16'b0011011011110111: color_data = 12'b001110100111;
		16'b0011011011111000: color_data = 12'b001110100111;
		16'b0011011011111001: color_data = 12'b001110100111;
		16'b0011011011111010: color_data = 12'b001110100111;
		16'b0011011011111011: color_data = 12'b001110100111;
		16'b0011011011111100: color_data = 12'b001110100111;
		16'b0011011011111101: color_data = 12'b001110100111;
		16'b0011011011111110: color_data = 12'b001110100111;
		16'b0011011011111111: color_data = 12'b001110100111;
		16'b0011011100000000: color_data = 12'b001110100111;
		16'b0011011100000001: color_data = 12'b001110100111;
		16'b0011011100011010: color_data = 12'b001110100111;
		16'b0011011100011011: color_data = 12'b001110100111;
		16'b0011011100011100: color_data = 12'b001110100111;
		16'b0011011100011101: color_data = 12'b001110100111;
		16'b0011011100011110: color_data = 12'b001110100111;
		16'b0011011100011111: color_data = 12'b001110100111;
		16'b0011011100100000: color_data = 12'b001110100111;
		16'b0011011100100001: color_data = 12'b001110100111;
		16'b0011011100100010: color_data = 12'b001110100111;
		16'b0011011100100011: color_data = 12'b001110100111;
		16'b0011011100100100: color_data = 12'b001110100111;
		16'b0011011100100101: color_data = 12'b001110100111;
		16'b0011011100100110: color_data = 12'b001110100111;
		16'b0011011100101101: color_data = 12'b001110100111;
		16'b0011011100101110: color_data = 12'b001110100111;
		16'b0011011100101111: color_data = 12'b001110100111;
		16'b0011011100110000: color_data = 12'b001110100111;
		16'b0011011100110001: color_data = 12'b001110100111;
		16'b0011011100110010: color_data = 12'b001110100111;
		16'b0011011100110011: color_data = 12'b001110100111;
		16'b0011011100110100: color_data = 12'b001110100111;
		16'b0011011100110101: color_data = 12'b001110100111;
		16'b0011011100110110: color_data = 12'b001110100111;
		16'b0011011100110111: color_data = 12'b001110100111;
		16'b0011011100111000: color_data = 12'b001110100111;
		16'b0011011101000101: color_data = 12'b001110100111;
		16'b0011011101000110: color_data = 12'b001110100111;
		16'b0011011101000111: color_data = 12'b001110100111;
		16'b0011011101001000: color_data = 12'b001110100111;
		16'b0011011101001001: color_data = 12'b001110100111;
		16'b0011011101001010: color_data = 12'b001110100111;
		16'b0011011101001011: color_data = 12'b001110100111;
		16'b0011011101001100: color_data = 12'b001110100111;
		16'b0011011101001101: color_data = 12'b001110100111;
		16'b0011011101001110: color_data = 12'b001110100111;
		16'b0011011101001111: color_data = 12'b001110100111;
		16'b0011011101010000: color_data = 12'b001110100111;
		16'b0011011101010001: color_data = 12'b001110100111;
		16'b0011011101011000: color_data = 12'b001110100111;
		16'b0011011101011001: color_data = 12'b001110100111;
		16'b0011011101011010: color_data = 12'b001110100111;
		16'b0011011101011011: color_data = 12'b001110100111;
		16'b0011011101011100: color_data = 12'b001110100111;
		16'b0011011101011101: color_data = 12'b001110100111;
		16'b0011011101011110: color_data = 12'b001110100111;
		16'b0011011101011111: color_data = 12'b001110100111;
		16'b0011011101100000: color_data = 12'b001110100111;
		16'b0011011101100001: color_data = 12'b001110100111;
		16'b0011011101100010: color_data = 12'b001110100111;
		16'b0011011101100011: color_data = 12'b001110100111;
		16'b0011100000000000: color_data = 12'b001110100111;
		16'b0011100000000001: color_data = 12'b001110100111;
		16'b0011100000000010: color_data = 12'b001110100111;
		16'b0011100000000011: color_data = 12'b001110100111;
		16'b0011100000000100: color_data = 12'b001110100111;
		16'b0011100000000101: color_data = 12'b001110100111;
		16'b0011100000000110: color_data = 12'b001110100111;
		16'b0011100000000111: color_data = 12'b001110100111;
		16'b0011100000001000: color_data = 12'b001110100111;
		16'b0011100000001001: color_data = 12'b001110100111;
		16'b0011100000001010: color_data = 12'b001110100111;
		16'b0011100000001011: color_data = 12'b001110100111;
		16'b0011100000001100: color_data = 12'b001110100111;
		16'b0011100000001101: color_data = 12'b001110100111;
		16'b0011100000001110: color_data = 12'b001110100111;
		16'b0011100000001111: color_data = 12'b001110100111;
		16'b0011100000010000: color_data = 12'b001110100111;
		16'b0011100000010001: color_data = 12'b001110100111;
		16'b0011100000010010: color_data = 12'b001110100111;
		16'b0011100000101011: color_data = 12'b001110100111;
		16'b0011100000101100: color_data = 12'b001110100111;
		16'b0011100000101101: color_data = 12'b001110100111;
		16'b0011100000101110: color_data = 12'b001110100111;
		16'b0011100000101111: color_data = 12'b001110100111;
		16'b0011100000110000: color_data = 12'b001110100111;
		16'b0011100000110001: color_data = 12'b001110100111;
		16'b0011100000110010: color_data = 12'b001110100111;
		16'b0011100000110011: color_data = 12'b001110100111;
		16'b0011100000110100: color_data = 12'b001110100111;
		16'b0011100000110101: color_data = 12'b001110100111;
		16'b0011100000110110: color_data = 12'b001110100111;
		16'b0011100000110111: color_data = 12'b001110100111;
		16'b0011100001000100: color_data = 12'b001110100111;
		16'b0011100001000101: color_data = 12'b001110100111;
		16'b0011100001000110: color_data = 12'b001110100111;
		16'b0011100001000111: color_data = 12'b001110100111;
		16'b0011100001001000: color_data = 12'b001110100111;
		16'b0011100001001001: color_data = 12'b001110100111;
		16'b0011100001001010: color_data = 12'b001110100111;
		16'b0011100001001011: color_data = 12'b001110100111;
		16'b0011100001001100: color_data = 12'b001110100111;
		16'b0011100001001101: color_data = 12'b001110100111;
		16'b0011100001001110: color_data = 12'b001110100111;
		16'b0011100001001111: color_data = 12'b001110100111;
		16'b0011100001011100: color_data = 12'b001110100111;
		16'b0011100001011101: color_data = 12'b001110100111;
		16'b0011100001011110: color_data = 12'b001110100111;
		16'b0011100001011111: color_data = 12'b001110100111;
		16'b0011100001100000: color_data = 12'b001110100111;
		16'b0011100001100001: color_data = 12'b001110100111;
		16'b0011100001100010: color_data = 12'b001110100111;
		16'b0011100001100011: color_data = 12'b001110100111;
		16'b0011100001100100: color_data = 12'b001110100111;
		16'b0011100001100101: color_data = 12'b001110100111;
		16'b0011100001100110: color_data = 12'b001110100111;
		16'b0011100001100111: color_data = 12'b001110100111;
		16'b0011100001101000: color_data = 12'b001110100111;
		16'b0011100001110101: color_data = 12'b001110100111;
		16'b0011100001110110: color_data = 12'b001110100111;
		16'b0011100001110111: color_data = 12'b001110100111;
		16'b0011100001111000: color_data = 12'b001110100111;
		16'b0011100001111001: color_data = 12'b001110100111;
		16'b0011100001111010: color_data = 12'b001110100111;
		16'b0011100001111011: color_data = 12'b001110100111;
		16'b0011100001111100: color_data = 12'b001110100111;
		16'b0011100001111101: color_data = 12'b001110100111;
		16'b0011100001111110: color_data = 12'b001110100111;
		16'b0011100001111111: color_data = 12'b001110100111;
		16'b0011100010000000: color_data = 12'b001110100111;
		16'b0011100010001101: color_data = 12'b001110100111;
		16'b0011100010001110: color_data = 12'b001110100111;
		16'b0011100010001111: color_data = 12'b001110100111;
		16'b0011100010010000: color_data = 12'b001110100111;
		16'b0011100010010001: color_data = 12'b001110100111;
		16'b0011100010010010: color_data = 12'b001110100111;
		16'b0011100010010011: color_data = 12'b001110100111;
		16'b0011100010010100: color_data = 12'b001110100111;
		16'b0011100010010101: color_data = 12'b001110100111;
		16'b0011100010010110: color_data = 12'b001110100111;
		16'b0011100010010111: color_data = 12'b001110100111;
		16'b0011100010011000: color_data = 12'b001110100111;
		16'b0011100010011001: color_data = 12'b001110100111;
		16'b0011100010100000: color_data = 12'b001110100111;
		16'b0011100010100001: color_data = 12'b001110100111;
		16'b0011100010100010: color_data = 12'b001110100111;
		16'b0011100010100011: color_data = 12'b001110100111;
		16'b0011100010100100: color_data = 12'b001110100111;
		16'b0011100010100101: color_data = 12'b001110100111;
		16'b0011100010100110: color_data = 12'b001110100111;
		16'b0011100010100111: color_data = 12'b001110100111;
		16'b0011100010101000: color_data = 12'b001110100111;
		16'b0011100010101001: color_data = 12'b001110100111;
		16'b0011100010101010: color_data = 12'b001110100111;
		16'b0011100010101011: color_data = 12'b001110100111;
		16'b0011100011001011: color_data = 12'b001110100111;
		16'b0011100011001100: color_data = 12'b001110100111;
		16'b0011100011001101: color_data = 12'b001110100111;
		16'b0011100011001110: color_data = 12'b001110100111;
		16'b0011100011001111: color_data = 12'b001110100111;
		16'b0011100011010000: color_data = 12'b001110100111;
		16'b0011100011010001: color_data = 12'b001110100111;
		16'b0011100011010010: color_data = 12'b001110100111;
		16'b0011100011010011: color_data = 12'b001110100111;
		16'b0011100011010100: color_data = 12'b001110100111;
		16'b0011100011010101: color_data = 12'b001110100111;
		16'b0011100011010110: color_data = 12'b001110100111;
		16'b0011100011100011: color_data = 12'b001110100111;
		16'b0011100011100100: color_data = 12'b001110100111;
		16'b0011100011100101: color_data = 12'b001110100111;
		16'b0011100011100110: color_data = 12'b001110100111;
		16'b0011100011100111: color_data = 12'b001110100111;
		16'b0011100011101000: color_data = 12'b001110100111;
		16'b0011100011101001: color_data = 12'b001110100111;
		16'b0011100011101010: color_data = 12'b001110100111;
		16'b0011100011101011: color_data = 12'b001110100111;
		16'b0011100011101100: color_data = 12'b001110100111;
		16'b0011100011101101: color_data = 12'b001110100111;
		16'b0011100011101110: color_data = 12'b001110100111;
		16'b0011100011101111: color_data = 12'b001110100111;
		16'b0011100011110110: color_data = 12'b001110100111;
		16'b0011100011110111: color_data = 12'b001110100111;
		16'b0011100011111000: color_data = 12'b001110100111;
		16'b0011100011111001: color_data = 12'b001110100111;
		16'b0011100011111010: color_data = 12'b001110100111;
		16'b0011100011111011: color_data = 12'b001110100111;
		16'b0011100011111100: color_data = 12'b001110100111;
		16'b0011100011111101: color_data = 12'b001110100111;
		16'b0011100011111110: color_data = 12'b001110100111;
		16'b0011100011111111: color_data = 12'b001110100111;
		16'b0011100100000000: color_data = 12'b001110100111;
		16'b0011100100000001: color_data = 12'b001110100111;
		16'b0011100100011010: color_data = 12'b001110100111;
		16'b0011100100011011: color_data = 12'b001110100111;
		16'b0011100100011100: color_data = 12'b001110100111;
		16'b0011100100011101: color_data = 12'b001110100111;
		16'b0011100100011110: color_data = 12'b001110100111;
		16'b0011100100011111: color_data = 12'b001110100111;
		16'b0011100100100000: color_data = 12'b001110100111;
		16'b0011100100100001: color_data = 12'b001110100111;
		16'b0011100100100010: color_data = 12'b001110100111;
		16'b0011100100100011: color_data = 12'b001110100111;
		16'b0011100100100100: color_data = 12'b001110100111;
		16'b0011100100100101: color_data = 12'b001110100111;
		16'b0011100100100110: color_data = 12'b001110100111;
		16'b0011100100101101: color_data = 12'b001110100111;
		16'b0011100100101110: color_data = 12'b001110100111;
		16'b0011100100101111: color_data = 12'b001110100111;
		16'b0011100100110000: color_data = 12'b001110100111;
		16'b0011100100110001: color_data = 12'b001110100111;
		16'b0011100100110010: color_data = 12'b001110100111;
		16'b0011100100110011: color_data = 12'b001110100111;
		16'b0011100100110100: color_data = 12'b001110100111;
		16'b0011100100110101: color_data = 12'b001110100111;
		16'b0011100100110110: color_data = 12'b001110100111;
		16'b0011100100110111: color_data = 12'b001110100111;
		16'b0011100100111000: color_data = 12'b001110100111;
		16'b0011100101000101: color_data = 12'b001110100111;
		16'b0011100101000110: color_data = 12'b001110100111;
		16'b0011100101000111: color_data = 12'b001110100111;
		16'b0011100101001000: color_data = 12'b001110100111;
		16'b0011100101001001: color_data = 12'b001110100111;
		16'b0011100101001010: color_data = 12'b001110100111;
		16'b0011100101001011: color_data = 12'b001110100111;
		16'b0011100101001100: color_data = 12'b001110100111;
		16'b0011100101001101: color_data = 12'b001110100111;
		16'b0011100101001110: color_data = 12'b001110100111;
		16'b0011100101001111: color_data = 12'b001110100111;
		16'b0011100101010000: color_data = 12'b001110100111;
		16'b0011100101010001: color_data = 12'b001110100111;
		16'b0011100101011000: color_data = 12'b001110100111;
		16'b0011100101011001: color_data = 12'b001110100111;
		16'b0011100101011010: color_data = 12'b001110100111;
		16'b0011100101011011: color_data = 12'b001110100111;
		16'b0011100101011100: color_data = 12'b001110100111;
		16'b0011100101011101: color_data = 12'b001110100111;
		16'b0011100101011110: color_data = 12'b001110100111;
		16'b0011100101011111: color_data = 12'b001110100111;
		16'b0011100101100000: color_data = 12'b001110100111;
		16'b0011100101100001: color_data = 12'b001110100111;
		16'b0011100101100010: color_data = 12'b001110100111;
		16'b0011100101100011: color_data = 12'b001110100111;
		16'b0011101000000000: color_data = 12'b001110100111;
		16'b0011101000000001: color_data = 12'b001110100111;
		16'b0011101000000010: color_data = 12'b001110100111;
		16'b0011101000000011: color_data = 12'b001110100111;
		16'b0011101000000100: color_data = 12'b001110100111;
		16'b0011101000000101: color_data = 12'b001110100111;
		16'b0011101000000110: color_data = 12'b001110100111;
		16'b0011101000000111: color_data = 12'b001110100111;
		16'b0011101000001000: color_data = 12'b001110100111;
		16'b0011101000001001: color_data = 12'b001110100111;
		16'b0011101000001010: color_data = 12'b001110100111;
		16'b0011101000001011: color_data = 12'b001110100111;
		16'b0011101000001100: color_data = 12'b001110100111;
		16'b0011101000001101: color_data = 12'b001110100111;
		16'b0011101000001110: color_data = 12'b001110100111;
		16'b0011101000001111: color_data = 12'b001110100111;
		16'b0011101000010000: color_data = 12'b001110100111;
		16'b0011101000010001: color_data = 12'b001110100111;
		16'b0011101000010010: color_data = 12'b001110100111;
		16'b0011101000101011: color_data = 12'b001110100111;
		16'b0011101000101100: color_data = 12'b001110100111;
		16'b0011101000101101: color_data = 12'b001110100111;
		16'b0011101000101110: color_data = 12'b001110100111;
		16'b0011101000101111: color_data = 12'b001110100111;
		16'b0011101000110000: color_data = 12'b001110100111;
		16'b0011101000110001: color_data = 12'b001110100111;
		16'b0011101000110010: color_data = 12'b001110100111;
		16'b0011101000110011: color_data = 12'b001110100111;
		16'b0011101000110100: color_data = 12'b001110100111;
		16'b0011101000110101: color_data = 12'b001110100111;
		16'b0011101000110110: color_data = 12'b001110100111;
		16'b0011101000110111: color_data = 12'b001110100111;
		16'b0011101001000100: color_data = 12'b001110100111;
		16'b0011101001000101: color_data = 12'b001110100111;
		16'b0011101001000110: color_data = 12'b001110100111;
		16'b0011101001000111: color_data = 12'b001110100111;
		16'b0011101001001000: color_data = 12'b001110100111;
		16'b0011101001001001: color_data = 12'b001110100111;
		16'b0011101001001010: color_data = 12'b001110100111;
		16'b0011101001001011: color_data = 12'b001110100111;
		16'b0011101001001100: color_data = 12'b001110100111;
		16'b0011101001001101: color_data = 12'b001110100111;
		16'b0011101001001110: color_data = 12'b001110100111;
		16'b0011101001001111: color_data = 12'b001110100111;
		16'b0011101001011100: color_data = 12'b001110100111;
		16'b0011101001011101: color_data = 12'b001110100111;
		16'b0011101001011110: color_data = 12'b001110100111;
		16'b0011101001011111: color_data = 12'b001110100111;
		16'b0011101001100000: color_data = 12'b001110100111;
		16'b0011101001100001: color_data = 12'b001110100111;
		16'b0011101001100010: color_data = 12'b001110100111;
		16'b0011101001100011: color_data = 12'b001110100111;
		16'b0011101001100100: color_data = 12'b001110100111;
		16'b0011101001100101: color_data = 12'b001110100111;
		16'b0011101001100110: color_data = 12'b001110100111;
		16'b0011101001100111: color_data = 12'b001110100111;
		16'b0011101001101000: color_data = 12'b001110100111;
		16'b0011101001110101: color_data = 12'b001110100111;
		16'b0011101001110110: color_data = 12'b001110100111;
		16'b0011101001110111: color_data = 12'b001110100111;
		16'b0011101001111000: color_data = 12'b001110100111;
		16'b0011101001111001: color_data = 12'b001110100111;
		16'b0011101001111010: color_data = 12'b001110100111;
		16'b0011101001111011: color_data = 12'b001110100111;
		16'b0011101001111100: color_data = 12'b001110100111;
		16'b0011101001111101: color_data = 12'b001110100111;
		16'b0011101001111110: color_data = 12'b001110100111;
		16'b0011101001111111: color_data = 12'b001110100111;
		16'b0011101010000000: color_data = 12'b001110100111;
		16'b0011101010001101: color_data = 12'b001110100111;
		16'b0011101010001110: color_data = 12'b001110100111;
		16'b0011101010001111: color_data = 12'b001110100111;
		16'b0011101010010000: color_data = 12'b001110100111;
		16'b0011101010010001: color_data = 12'b001110100111;
		16'b0011101010010010: color_data = 12'b001110100111;
		16'b0011101010010011: color_data = 12'b001110100111;
		16'b0011101010010100: color_data = 12'b001110100111;
		16'b0011101010010101: color_data = 12'b001110100111;
		16'b0011101010010110: color_data = 12'b001110100111;
		16'b0011101010010111: color_data = 12'b001110100111;
		16'b0011101010011000: color_data = 12'b001110100111;
		16'b0011101010011001: color_data = 12'b001110100111;
		16'b0011101010100000: color_data = 12'b001110100111;
		16'b0011101010100001: color_data = 12'b001110100111;
		16'b0011101010100010: color_data = 12'b001110100111;
		16'b0011101010100011: color_data = 12'b001110100111;
		16'b0011101010100100: color_data = 12'b001110100111;
		16'b0011101010100101: color_data = 12'b001110100111;
		16'b0011101010100110: color_data = 12'b001110100111;
		16'b0011101010100111: color_data = 12'b001110100111;
		16'b0011101010101000: color_data = 12'b001110100111;
		16'b0011101010101001: color_data = 12'b001110100111;
		16'b0011101010101010: color_data = 12'b001110100111;
		16'b0011101010101011: color_data = 12'b001110100111;
		16'b0011101011001011: color_data = 12'b001110100111;
		16'b0011101011001100: color_data = 12'b001110100111;
		16'b0011101011001101: color_data = 12'b001110100111;
		16'b0011101011001110: color_data = 12'b001110100111;
		16'b0011101011001111: color_data = 12'b001110100111;
		16'b0011101011010000: color_data = 12'b001110100111;
		16'b0011101011010001: color_data = 12'b001110100111;
		16'b0011101011010010: color_data = 12'b001110100111;
		16'b0011101011010011: color_data = 12'b001110100111;
		16'b0011101011010100: color_data = 12'b001110100111;
		16'b0011101011010101: color_data = 12'b001110100111;
		16'b0011101011010110: color_data = 12'b001110100111;
		16'b0011101011100011: color_data = 12'b001110100111;
		16'b0011101011100100: color_data = 12'b001110100111;
		16'b0011101011100101: color_data = 12'b001110100111;
		16'b0011101011100110: color_data = 12'b001110100111;
		16'b0011101011100111: color_data = 12'b001110100111;
		16'b0011101011101000: color_data = 12'b001110100111;
		16'b0011101011101001: color_data = 12'b001110100111;
		16'b0011101011101010: color_data = 12'b001110100111;
		16'b0011101011101011: color_data = 12'b001110100111;
		16'b0011101011101100: color_data = 12'b001110100111;
		16'b0011101011101101: color_data = 12'b001110100111;
		16'b0011101011101110: color_data = 12'b001110100111;
		16'b0011101011101111: color_data = 12'b001110100111;
		16'b0011101011110110: color_data = 12'b001110100111;
		16'b0011101011110111: color_data = 12'b001110100111;
		16'b0011101011111000: color_data = 12'b001110100111;
		16'b0011101011111001: color_data = 12'b001110100111;
		16'b0011101011111010: color_data = 12'b001110100111;
		16'b0011101011111011: color_data = 12'b001110100111;
		16'b0011101011111100: color_data = 12'b001110100111;
		16'b0011101011111101: color_data = 12'b001110100111;
		16'b0011101011111110: color_data = 12'b001110100111;
		16'b0011101011111111: color_data = 12'b001110100111;
		16'b0011101100000000: color_data = 12'b001110100111;
		16'b0011101100000001: color_data = 12'b001110100111;
		16'b0011101100011010: color_data = 12'b001110100111;
		16'b0011101100011011: color_data = 12'b001110100111;
		16'b0011101100011100: color_data = 12'b001110100111;
		16'b0011101100011101: color_data = 12'b001110100111;
		16'b0011101100011110: color_data = 12'b001110100111;
		16'b0011101100011111: color_data = 12'b001110100111;
		16'b0011101100100000: color_data = 12'b001110100111;
		16'b0011101100100001: color_data = 12'b001110100111;
		16'b0011101100100010: color_data = 12'b001110100111;
		16'b0011101100100011: color_data = 12'b001110100111;
		16'b0011101100100100: color_data = 12'b001110100111;
		16'b0011101100100101: color_data = 12'b001110100111;
		16'b0011101100100110: color_data = 12'b001110100111;
		16'b0011101100101101: color_data = 12'b001110100111;
		16'b0011101100101110: color_data = 12'b001110100111;
		16'b0011101100101111: color_data = 12'b001110100111;
		16'b0011101100110000: color_data = 12'b001110100111;
		16'b0011101100110001: color_data = 12'b001110100111;
		16'b0011101100110010: color_data = 12'b001110100111;
		16'b0011101100110011: color_data = 12'b001110100111;
		16'b0011101100110100: color_data = 12'b001110100111;
		16'b0011101100110101: color_data = 12'b001110100111;
		16'b0011101100110110: color_data = 12'b001110100111;
		16'b0011101100110111: color_data = 12'b001110100111;
		16'b0011101100111000: color_data = 12'b001110100111;
		16'b0011101101000101: color_data = 12'b001110100111;
		16'b0011101101000110: color_data = 12'b001110100111;
		16'b0011101101000111: color_data = 12'b001110100111;
		16'b0011101101001000: color_data = 12'b001110100111;
		16'b0011101101001001: color_data = 12'b001110100111;
		16'b0011101101001010: color_data = 12'b001110100111;
		16'b0011101101001011: color_data = 12'b001110100111;
		16'b0011101101001100: color_data = 12'b001110100111;
		16'b0011101101001101: color_data = 12'b001110100111;
		16'b0011101101001110: color_data = 12'b001110100111;
		16'b0011101101001111: color_data = 12'b001110100111;
		16'b0011101101010000: color_data = 12'b001110100111;
		16'b0011101101010001: color_data = 12'b001110100111;
		16'b0011101101011000: color_data = 12'b001110100111;
		16'b0011101101011001: color_data = 12'b001110100111;
		16'b0011101101011010: color_data = 12'b001110100111;
		16'b0011101101011011: color_data = 12'b001110100111;
		16'b0011101101011100: color_data = 12'b001110100111;
		16'b0011101101011101: color_data = 12'b001110100111;
		16'b0011101101011110: color_data = 12'b001110100111;
		16'b0011101101011111: color_data = 12'b001110100111;
		16'b0011101101100000: color_data = 12'b001110100111;
		16'b0011101101100001: color_data = 12'b001110100111;
		16'b0011101101100010: color_data = 12'b001110100111;
		16'b0011101101100011: color_data = 12'b001110100111;
		16'b0011110000000000: color_data = 12'b001110100111;
		16'b0011110000000001: color_data = 12'b001110100111;
		16'b0011110000000010: color_data = 12'b001110100111;
		16'b0011110000000011: color_data = 12'b001110100111;
		16'b0011110000000100: color_data = 12'b001110100111;
		16'b0011110000000101: color_data = 12'b001110100111;
		16'b0011110000000110: color_data = 12'b001110100111;
		16'b0011110000000111: color_data = 12'b001110100111;
		16'b0011110000001000: color_data = 12'b001110100111;
		16'b0011110000001001: color_data = 12'b001110100111;
		16'b0011110000001010: color_data = 12'b001110100111;
		16'b0011110000001011: color_data = 12'b001110100111;
		16'b0011110000001100: color_data = 12'b001110100111;
		16'b0011110000001101: color_data = 12'b001110100111;
		16'b0011110000001110: color_data = 12'b001110100111;
		16'b0011110000001111: color_data = 12'b001110100111;
		16'b0011110000010000: color_data = 12'b001110100111;
		16'b0011110000010001: color_data = 12'b001110100111;
		16'b0011110000010010: color_data = 12'b001110100111;
		16'b0011110000101011: color_data = 12'b001110100111;
		16'b0011110000101100: color_data = 12'b001110100111;
		16'b0011110000101101: color_data = 12'b001110100111;
		16'b0011110000101110: color_data = 12'b001110100111;
		16'b0011110000101111: color_data = 12'b001110100111;
		16'b0011110000110000: color_data = 12'b001110100111;
		16'b0011110000110001: color_data = 12'b001110100111;
		16'b0011110000110010: color_data = 12'b001110100111;
		16'b0011110000110011: color_data = 12'b001110100111;
		16'b0011110000110100: color_data = 12'b001110100111;
		16'b0011110000110101: color_data = 12'b001110100111;
		16'b0011110000110110: color_data = 12'b001110100111;
		16'b0011110000110111: color_data = 12'b001110100111;
		16'b0011110001000100: color_data = 12'b001110100111;
		16'b0011110001000101: color_data = 12'b001110100111;
		16'b0011110001000110: color_data = 12'b001110100111;
		16'b0011110001000111: color_data = 12'b001110100111;
		16'b0011110001001000: color_data = 12'b001110100111;
		16'b0011110001001001: color_data = 12'b001110100111;
		16'b0011110001001010: color_data = 12'b001110100111;
		16'b0011110001001011: color_data = 12'b001110100111;
		16'b0011110001001100: color_data = 12'b001110100111;
		16'b0011110001001101: color_data = 12'b001110100111;
		16'b0011110001001110: color_data = 12'b001110100111;
		16'b0011110001001111: color_data = 12'b001110100111;
		16'b0011110001011100: color_data = 12'b001110100111;
		16'b0011110001011101: color_data = 12'b001110100111;
		16'b0011110001011110: color_data = 12'b001110100111;
		16'b0011110001011111: color_data = 12'b001110100111;
		16'b0011110001100000: color_data = 12'b001110100111;
		16'b0011110001100001: color_data = 12'b001110100111;
		16'b0011110001100010: color_data = 12'b001110100111;
		16'b0011110001100011: color_data = 12'b001110100111;
		16'b0011110001100100: color_data = 12'b001110100111;
		16'b0011110001100101: color_data = 12'b001110100111;
		16'b0011110001100110: color_data = 12'b001110100111;
		16'b0011110001100111: color_data = 12'b001110100111;
		16'b0011110001101000: color_data = 12'b001110100111;
		16'b0011110001110101: color_data = 12'b001110100111;
		16'b0011110001110110: color_data = 12'b001110100111;
		16'b0011110001110111: color_data = 12'b001110100111;
		16'b0011110001111000: color_data = 12'b001110100111;
		16'b0011110001111001: color_data = 12'b001110100111;
		16'b0011110001111010: color_data = 12'b001110100111;
		16'b0011110001111011: color_data = 12'b001110100111;
		16'b0011110001111100: color_data = 12'b001110100111;
		16'b0011110001111101: color_data = 12'b001110100111;
		16'b0011110001111110: color_data = 12'b001110100111;
		16'b0011110001111111: color_data = 12'b001110100111;
		16'b0011110010000000: color_data = 12'b001110100111;
		16'b0011110010001101: color_data = 12'b001110100111;
		16'b0011110010001110: color_data = 12'b001110100111;
		16'b0011110010001111: color_data = 12'b001110100111;
		16'b0011110010010000: color_data = 12'b001110100111;
		16'b0011110010010001: color_data = 12'b001110100111;
		16'b0011110010010010: color_data = 12'b001110100111;
		16'b0011110010010011: color_data = 12'b001110100111;
		16'b0011110010010100: color_data = 12'b001110100111;
		16'b0011110010010101: color_data = 12'b001110100111;
		16'b0011110010010110: color_data = 12'b001110100111;
		16'b0011110010010111: color_data = 12'b001110100111;
		16'b0011110010011000: color_data = 12'b001110100111;
		16'b0011110010011001: color_data = 12'b001110100111;
		16'b0011110010100000: color_data = 12'b001110100111;
		16'b0011110010100001: color_data = 12'b001110100111;
		16'b0011110010100010: color_data = 12'b001110100111;
		16'b0011110010100011: color_data = 12'b001110100111;
		16'b0011110010100100: color_data = 12'b001110100111;
		16'b0011110010100101: color_data = 12'b001110100111;
		16'b0011110010100110: color_data = 12'b001110100111;
		16'b0011110010100111: color_data = 12'b001110100111;
		16'b0011110010101000: color_data = 12'b001110100111;
		16'b0011110010101001: color_data = 12'b001110100111;
		16'b0011110010101010: color_data = 12'b001110100111;
		16'b0011110010101011: color_data = 12'b001110100111;
		16'b0011110011001011: color_data = 12'b001110100111;
		16'b0011110011001100: color_data = 12'b001110100111;
		16'b0011110011001101: color_data = 12'b001110100111;
		16'b0011110011001110: color_data = 12'b001110100111;
		16'b0011110011001111: color_data = 12'b001110100111;
		16'b0011110011010000: color_data = 12'b001110100111;
		16'b0011110011010001: color_data = 12'b001110100111;
		16'b0011110011010010: color_data = 12'b001110100111;
		16'b0011110011010011: color_data = 12'b001110100111;
		16'b0011110011010100: color_data = 12'b001110100111;
		16'b0011110011010101: color_data = 12'b001110100111;
		16'b0011110011010110: color_data = 12'b001110100111;
		16'b0011110011100011: color_data = 12'b001110100111;
		16'b0011110011100100: color_data = 12'b001110100111;
		16'b0011110011100101: color_data = 12'b001110100111;
		16'b0011110011100110: color_data = 12'b001110100111;
		16'b0011110011100111: color_data = 12'b001110100111;
		16'b0011110011101000: color_data = 12'b001110100111;
		16'b0011110011101001: color_data = 12'b001110100111;
		16'b0011110011101010: color_data = 12'b001110100111;
		16'b0011110011101011: color_data = 12'b001110100111;
		16'b0011110011101100: color_data = 12'b001110100111;
		16'b0011110011101101: color_data = 12'b001110100111;
		16'b0011110011101110: color_data = 12'b001110100111;
		16'b0011110011101111: color_data = 12'b001110100111;
		16'b0011110011110110: color_data = 12'b001110100111;
		16'b0011110011110111: color_data = 12'b001110100111;
		16'b0011110011111000: color_data = 12'b001110100111;
		16'b0011110011111001: color_data = 12'b001110100111;
		16'b0011110011111010: color_data = 12'b001110100111;
		16'b0011110011111011: color_data = 12'b001110100111;
		16'b0011110011111100: color_data = 12'b001110100111;
		16'b0011110011111101: color_data = 12'b001110100111;
		16'b0011110011111110: color_data = 12'b001110100111;
		16'b0011110011111111: color_data = 12'b001110100111;
		16'b0011110100000000: color_data = 12'b001110100111;
		16'b0011110100000001: color_data = 12'b001110100111;
		16'b0011110100011010: color_data = 12'b001110100111;
		16'b0011110100011011: color_data = 12'b001110100111;
		16'b0011110100011100: color_data = 12'b001110100111;
		16'b0011110100011101: color_data = 12'b001110100111;
		16'b0011110100011110: color_data = 12'b001110100111;
		16'b0011110100011111: color_data = 12'b001110100111;
		16'b0011110100100000: color_data = 12'b001110100111;
		16'b0011110100100001: color_data = 12'b001110100111;
		16'b0011110100100010: color_data = 12'b001110100111;
		16'b0011110100100011: color_data = 12'b001110100111;
		16'b0011110100100100: color_data = 12'b001110100111;
		16'b0011110100100101: color_data = 12'b001110100111;
		16'b0011110100100110: color_data = 12'b001110100111;
		16'b0011110100101101: color_data = 12'b001110100111;
		16'b0011110100101110: color_data = 12'b001110100111;
		16'b0011110100101111: color_data = 12'b001110100111;
		16'b0011110100110000: color_data = 12'b001110100111;
		16'b0011110100110001: color_data = 12'b001110100111;
		16'b0011110100110010: color_data = 12'b001110100111;
		16'b0011110100110011: color_data = 12'b001110100111;
		16'b0011110100110100: color_data = 12'b001110100111;
		16'b0011110100110101: color_data = 12'b001110100111;
		16'b0011110100110110: color_data = 12'b001110100111;
		16'b0011110100110111: color_data = 12'b001110100111;
		16'b0011110100111000: color_data = 12'b001110100111;
		16'b0011110101000101: color_data = 12'b001110100111;
		16'b0011110101000110: color_data = 12'b001110100111;
		16'b0011110101000111: color_data = 12'b001110100111;
		16'b0011110101001000: color_data = 12'b001110100111;
		16'b0011110101001001: color_data = 12'b001110100111;
		16'b0011110101001010: color_data = 12'b001110100111;
		16'b0011110101001011: color_data = 12'b001110100111;
		16'b0011110101001100: color_data = 12'b001110100111;
		16'b0011110101001101: color_data = 12'b001110100111;
		16'b0011110101001110: color_data = 12'b001110100111;
		16'b0011110101001111: color_data = 12'b001110100111;
		16'b0011110101010000: color_data = 12'b001110100111;
		16'b0011110101010001: color_data = 12'b001110100111;
		16'b0011110101011000: color_data = 12'b001110100111;
		16'b0011110101011001: color_data = 12'b001110100111;
		16'b0011110101011010: color_data = 12'b001110100111;
		16'b0011110101011011: color_data = 12'b001110100111;
		16'b0011110101011100: color_data = 12'b001110100111;
		16'b0011110101011101: color_data = 12'b001110100111;
		16'b0011110101011110: color_data = 12'b001110100111;
		16'b0011110101011111: color_data = 12'b001110100111;
		16'b0011110101100000: color_data = 12'b001110100111;
		16'b0011110101100001: color_data = 12'b001110100111;
		16'b0011110101100010: color_data = 12'b001110100111;
		16'b0011110101100011: color_data = 12'b001110100111;
		16'b0011111000000000: color_data = 12'b001110100111;
		16'b0011111000000001: color_data = 12'b001110100111;
		16'b0011111000000010: color_data = 12'b001110100111;
		16'b0011111000000011: color_data = 12'b001110100111;
		16'b0011111000000100: color_data = 12'b001110100111;
		16'b0011111000000101: color_data = 12'b001110100111;
		16'b0011111000000110: color_data = 12'b001110100111;
		16'b0011111000000111: color_data = 12'b001110100111;
		16'b0011111000001000: color_data = 12'b001110100111;
		16'b0011111000001001: color_data = 12'b001110100111;
		16'b0011111000001010: color_data = 12'b001110100111;
		16'b0011111000001011: color_data = 12'b001110100111;
		16'b0011111000001100: color_data = 12'b001110100111;
		16'b0011111000001101: color_data = 12'b001110100111;
		16'b0011111000001110: color_data = 12'b001110100111;
		16'b0011111000001111: color_data = 12'b001110100111;
		16'b0011111000010000: color_data = 12'b001110100111;
		16'b0011111000010001: color_data = 12'b001110100111;
		16'b0011111000010010: color_data = 12'b001110100111;
		16'b0011111000101011: color_data = 12'b001110100111;
		16'b0011111000101100: color_data = 12'b001110100111;
		16'b0011111000101101: color_data = 12'b001110100111;
		16'b0011111000101110: color_data = 12'b001110100111;
		16'b0011111000101111: color_data = 12'b001110100111;
		16'b0011111000110000: color_data = 12'b001110100111;
		16'b0011111000110001: color_data = 12'b001110100111;
		16'b0011111000110010: color_data = 12'b001110100111;
		16'b0011111000110011: color_data = 12'b001110100111;
		16'b0011111000110100: color_data = 12'b001110100111;
		16'b0011111000110101: color_data = 12'b001110100111;
		16'b0011111000110110: color_data = 12'b001110100111;
		16'b0011111000110111: color_data = 12'b001110100111;
		16'b0011111001000100: color_data = 12'b001110100111;
		16'b0011111001000101: color_data = 12'b001110100111;
		16'b0011111001000110: color_data = 12'b001110100111;
		16'b0011111001000111: color_data = 12'b001110100111;
		16'b0011111001001000: color_data = 12'b001110100111;
		16'b0011111001001001: color_data = 12'b001110100111;
		16'b0011111001001010: color_data = 12'b001110100111;
		16'b0011111001001011: color_data = 12'b001110100111;
		16'b0011111001001100: color_data = 12'b001110100111;
		16'b0011111001001101: color_data = 12'b001110100111;
		16'b0011111001001110: color_data = 12'b001110100111;
		16'b0011111001001111: color_data = 12'b001110100111;
		16'b0011111001011100: color_data = 12'b001110100111;
		16'b0011111001011101: color_data = 12'b001110100111;
		16'b0011111001011110: color_data = 12'b001110100111;
		16'b0011111001011111: color_data = 12'b001110100111;
		16'b0011111001100000: color_data = 12'b001110100111;
		16'b0011111001100001: color_data = 12'b001110100111;
		16'b0011111001100010: color_data = 12'b001110100111;
		16'b0011111001100011: color_data = 12'b001110100111;
		16'b0011111001100100: color_data = 12'b001110100111;
		16'b0011111001100101: color_data = 12'b001110100111;
		16'b0011111001100110: color_data = 12'b001110100111;
		16'b0011111001100111: color_data = 12'b001110100111;
		16'b0011111001101000: color_data = 12'b001110100111;
		16'b0011111001110101: color_data = 12'b001110100111;
		16'b0011111001110110: color_data = 12'b001110100111;
		16'b0011111001110111: color_data = 12'b001110100111;
		16'b0011111001111000: color_data = 12'b001110100111;
		16'b0011111001111001: color_data = 12'b001110100111;
		16'b0011111001111010: color_data = 12'b001110100111;
		16'b0011111001111011: color_data = 12'b001110100111;
		16'b0011111001111100: color_data = 12'b001110100111;
		16'b0011111001111101: color_data = 12'b001110100111;
		16'b0011111001111110: color_data = 12'b001110100111;
		16'b0011111001111111: color_data = 12'b001110100111;
		16'b0011111010000000: color_data = 12'b001110100111;
		16'b0011111010001101: color_data = 12'b001110100111;
		16'b0011111010001110: color_data = 12'b001110100111;
		16'b0011111010001111: color_data = 12'b001110100111;
		16'b0011111010010000: color_data = 12'b001110100111;
		16'b0011111010010001: color_data = 12'b001110100111;
		16'b0011111010010010: color_data = 12'b001110100111;
		16'b0011111010010011: color_data = 12'b001110100111;
		16'b0011111010010100: color_data = 12'b001110100111;
		16'b0011111010010101: color_data = 12'b001110100111;
		16'b0011111010010110: color_data = 12'b001110100111;
		16'b0011111010010111: color_data = 12'b001110100111;
		16'b0011111010011000: color_data = 12'b001110100111;
		16'b0011111010011001: color_data = 12'b001110100111;
		16'b0011111010100000: color_data = 12'b001110100111;
		16'b0011111010100001: color_data = 12'b001110100111;
		16'b0011111010100010: color_data = 12'b001110100111;
		16'b0011111010100011: color_data = 12'b001110100111;
		16'b0011111010100100: color_data = 12'b001110100111;
		16'b0011111010100101: color_data = 12'b001110100111;
		16'b0011111010100110: color_data = 12'b001110100111;
		16'b0011111010100111: color_data = 12'b001110100111;
		16'b0011111010101000: color_data = 12'b001110100111;
		16'b0011111010101001: color_data = 12'b001110100111;
		16'b0011111010101010: color_data = 12'b001110100111;
		16'b0011111010101011: color_data = 12'b001110100111;
		16'b0011111011001011: color_data = 12'b001110100111;
		16'b0011111011001100: color_data = 12'b001110100111;
		16'b0011111011001101: color_data = 12'b001110100111;
		16'b0011111011001110: color_data = 12'b001110100111;
		16'b0011111011001111: color_data = 12'b001110100111;
		16'b0011111011010000: color_data = 12'b001110100111;
		16'b0011111011010001: color_data = 12'b001110100111;
		16'b0011111011010010: color_data = 12'b001110100111;
		16'b0011111011010011: color_data = 12'b001110100111;
		16'b0011111011010100: color_data = 12'b001110100111;
		16'b0011111011010101: color_data = 12'b001110100111;
		16'b0011111011010110: color_data = 12'b001110100111;
		16'b0011111011100011: color_data = 12'b001110100111;
		16'b0011111011100100: color_data = 12'b001110100111;
		16'b0011111011100101: color_data = 12'b001110100111;
		16'b0011111011100110: color_data = 12'b001110100111;
		16'b0011111011100111: color_data = 12'b001110100111;
		16'b0011111011101000: color_data = 12'b001110100111;
		16'b0011111011101001: color_data = 12'b001110100111;
		16'b0011111011101010: color_data = 12'b001110100111;
		16'b0011111011101011: color_data = 12'b001110100111;
		16'b0011111011101100: color_data = 12'b001110100111;
		16'b0011111011101101: color_data = 12'b001110100111;
		16'b0011111011101110: color_data = 12'b001110100111;
		16'b0011111011101111: color_data = 12'b001110100111;
		16'b0011111011110110: color_data = 12'b001110100111;
		16'b0011111011110111: color_data = 12'b001110100111;
		16'b0011111011111000: color_data = 12'b001110100111;
		16'b0011111011111001: color_data = 12'b001110100111;
		16'b0011111011111010: color_data = 12'b001110100111;
		16'b0011111011111011: color_data = 12'b001110100111;
		16'b0011111011111100: color_data = 12'b001110100111;
		16'b0011111011111101: color_data = 12'b001110100111;
		16'b0011111011111110: color_data = 12'b001110100111;
		16'b0011111011111111: color_data = 12'b001110100111;
		16'b0011111100000000: color_data = 12'b001110100111;
		16'b0011111100000001: color_data = 12'b001110100111;
		16'b0011111100011010: color_data = 12'b001110100111;
		16'b0011111100011011: color_data = 12'b001110100111;
		16'b0011111100011100: color_data = 12'b001110100111;
		16'b0011111100011101: color_data = 12'b001110100111;
		16'b0011111100011110: color_data = 12'b001110100111;
		16'b0011111100011111: color_data = 12'b001110100111;
		16'b0011111100100000: color_data = 12'b001110100111;
		16'b0011111100100001: color_data = 12'b001110100111;
		16'b0011111100100010: color_data = 12'b001110100111;
		16'b0011111100100011: color_data = 12'b001110100111;
		16'b0011111100100100: color_data = 12'b001110100111;
		16'b0011111100100101: color_data = 12'b001110100111;
		16'b0011111100100110: color_data = 12'b001110100111;
		16'b0011111100101101: color_data = 12'b001110100111;
		16'b0011111100101110: color_data = 12'b001110100111;
		16'b0011111100101111: color_data = 12'b001110100111;
		16'b0011111100110000: color_data = 12'b001110100111;
		16'b0011111100110001: color_data = 12'b001110100111;
		16'b0011111100110010: color_data = 12'b001110100111;
		16'b0011111100110011: color_data = 12'b001110100111;
		16'b0011111100110100: color_data = 12'b001110100111;
		16'b0011111100110101: color_data = 12'b001110100111;
		16'b0011111100110110: color_data = 12'b001110100111;
		16'b0011111100110111: color_data = 12'b001110100111;
		16'b0011111100111000: color_data = 12'b001110100111;
		16'b0011111101000101: color_data = 12'b001110100111;
		16'b0011111101000110: color_data = 12'b001110100111;
		16'b0011111101000111: color_data = 12'b001110100111;
		16'b0011111101001000: color_data = 12'b001110100111;
		16'b0011111101001001: color_data = 12'b001110100111;
		16'b0011111101001010: color_data = 12'b001110100111;
		16'b0011111101001011: color_data = 12'b001110100111;
		16'b0011111101001100: color_data = 12'b001110100111;
		16'b0011111101001101: color_data = 12'b001110100111;
		16'b0011111101001110: color_data = 12'b001110100111;
		16'b0011111101001111: color_data = 12'b001110100111;
		16'b0011111101010000: color_data = 12'b001110100111;
		16'b0011111101010001: color_data = 12'b001110100111;
		16'b0011111101011000: color_data = 12'b001110100111;
		16'b0011111101011001: color_data = 12'b001110100111;
		16'b0011111101011010: color_data = 12'b001110100111;
		16'b0011111101011011: color_data = 12'b001110100111;
		16'b0011111101011100: color_data = 12'b001110100111;
		16'b0011111101011101: color_data = 12'b001110100111;
		16'b0011111101011110: color_data = 12'b001110100111;
		16'b0011111101011111: color_data = 12'b001110100111;
		16'b0011111101100000: color_data = 12'b001110100111;
		16'b0011111101100001: color_data = 12'b001110100111;
		16'b0011111101100010: color_data = 12'b001110100111;
		16'b0011111101100011: color_data = 12'b001110100111;
		16'b0100000000000000: color_data = 12'b001110100111;
		16'b0100000000000001: color_data = 12'b001110100111;
		16'b0100000000000010: color_data = 12'b001110100111;
		16'b0100000000000011: color_data = 12'b001110100111;
		16'b0100000000000100: color_data = 12'b001110100111;
		16'b0100000000000101: color_data = 12'b001110100111;
		16'b0100000000000110: color_data = 12'b001110100111;
		16'b0100000000000111: color_data = 12'b001110100111;
		16'b0100000000001000: color_data = 12'b001110100111;
		16'b0100000000001001: color_data = 12'b001110100111;
		16'b0100000000001010: color_data = 12'b001110100111;
		16'b0100000000001011: color_data = 12'b001110100111;
		16'b0100000000001100: color_data = 12'b001110100111;
		16'b0100000000001101: color_data = 12'b001110100111;
		16'b0100000000001110: color_data = 12'b001110100111;
		16'b0100000000001111: color_data = 12'b001110100111;
		16'b0100000000010000: color_data = 12'b001110100111;
		16'b0100000000010001: color_data = 12'b001110100111;
		16'b0100000000010010: color_data = 12'b001110100111;
		16'b0100000000101011: color_data = 12'b001110100111;
		16'b0100000000101100: color_data = 12'b001110100111;
		16'b0100000000101101: color_data = 12'b001110100111;
		16'b0100000000101110: color_data = 12'b001110100111;
		16'b0100000000101111: color_data = 12'b001110100111;
		16'b0100000000110000: color_data = 12'b001110100111;
		16'b0100000000110001: color_data = 12'b001110100111;
		16'b0100000000110010: color_data = 12'b001110100111;
		16'b0100000000110011: color_data = 12'b001110100111;
		16'b0100000000110100: color_data = 12'b001110100111;
		16'b0100000000110101: color_data = 12'b001110100111;
		16'b0100000000110110: color_data = 12'b001110100111;
		16'b0100000000110111: color_data = 12'b001110100111;
		16'b0100000001000100: color_data = 12'b001110100111;
		16'b0100000001000101: color_data = 12'b001110100111;
		16'b0100000001000110: color_data = 12'b001110100111;
		16'b0100000001000111: color_data = 12'b001110100111;
		16'b0100000001001000: color_data = 12'b001110100111;
		16'b0100000001001001: color_data = 12'b001110100111;
		16'b0100000001001010: color_data = 12'b001110100111;
		16'b0100000001001011: color_data = 12'b001110100111;
		16'b0100000001001100: color_data = 12'b001110100111;
		16'b0100000001001101: color_data = 12'b001110100111;
		16'b0100000001001110: color_data = 12'b001110100111;
		16'b0100000001001111: color_data = 12'b001110100111;
		16'b0100000001011100: color_data = 12'b001110100111;
		16'b0100000001011101: color_data = 12'b001110100111;
		16'b0100000001011110: color_data = 12'b001110100111;
		16'b0100000001011111: color_data = 12'b001110100111;
		16'b0100000001100000: color_data = 12'b001110100111;
		16'b0100000001100001: color_data = 12'b001110100111;
		16'b0100000001100010: color_data = 12'b001110100111;
		16'b0100000001100011: color_data = 12'b001110100111;
		16'b0100000001100100: color_data = 12'b001110100111;
		16'b0100000001100101: color_data = 12'b001110100111;
		16'b0100000001100110: color_data = 12'b001110100111;
		16'b0100000001100111: color_data = 12'b001110100111;
		16'b0100000001101000: color_data = 12'b001110100111;
		16'b0100000001110101: color_data = 12'b001110100111;
		16'b0100000001110110: color_data = 12'b001110100111;
		16'b0100000001110111: color_data = 12'b001110100111;
		16'b0100000001111000: color_data = 12'b001110100111;
		16'b0100000001111001: color_data = 12'b001110100111;
		16'b0100000001111010: color_data = 12'b001110100111;
		16'b0100000001111011: color_data = 12'b001110100111;
		16'b0100000001111100: color_data = 12'b001110100111;
		16'b0100000001111101: color_data = 12'b001110100111;
		16'b0100000001111110: color_data = 12'b001110100111;
		16'b0100000001111111: color_data = 12'b001110100111;
		16'b0100000010000000: color_data = 12'b001110100111;
		16'b0100000010001101: color_data = 12'b001110100111;
		16'b0100000010001110: color_data = 12'b001110100111;
		16'b0100000010001111: color_data = 12'b001110100111;
		16'b0100000010010000: color_data = 12'b001110100111;
		16'b0100000010010001: color_data = 12'b001110100111;
		16'b0100000010010010: color_data = 12'b001110100111;
		16'b0100000010010011: color_data = 12'b001110100111;
		16'b0100000010010100: color_data = 12'b001110100111;
		16'b0100000010010101: color_data = 12'b001110100111;
		16'b0100000010010110: color_data = 12'b001110100111;
		16'b0100000010010111: color_data = 12'b001110100111;
		16'b0100000010011000: color_data = 12'b001110100111;
		16'b0100000010011001: color_data = 12'b001110100111;
		16'b0100000010100000: color_data = 12'b001110100111;
		16'b0100000010100001: color_data = 12'b001110100111;
		16'b0100000010100010: color_data = 12'b001110100111;
		16'b0100000010100011: color_data = 12'b001110100111;
		16'b0100000010100100: color_data = 12'b001110100111;
		16'b0100000010100101: color_data = 12'b001110100111;
		16'b0100000010100110: color_data = 12'b001110100111;
		16'b0100000010100111: color_data = 12'b001110100111;
		16'b0100000010101000: color_data = 12'b001110100111;
		16'b0100000010101001: color_data = 12'b001110100111;
		16'b0100000010101010: color_data = 12'b001110100111;
		16'b0100000010101011: color_data = 12'b001110100111;
		16'b0100000011001011: color_data = 12'b001110100111;
		16'b0100000011001100: color_data = 12'b001110100111;
		16'b0100000011001101: color_data = 12'b001110100111;
		16'b0100000011001110: color_data = 12'b001110100111;
		16'b0100000011001111: color_data = 12'b001110100111;
		16'b0100000011010000: color_data = 12'b001110100111;
		16'b0100000011010001: color_data = 12'b001110100111;
		16'b0100000011010010: color_data = 12'b001110100111;
		16'b0100000011010011: color_data = 12'b001110100111;
		16'b0100000011010100: color_data = 12'b001110100111;
		16'b0100000011010101: color_data = 12'b001110100111;
		16'b0100000011010110: color_data = 12'b001110100111;
		16'b0100000011100011: color_data = 12'b001110100111;
		16'b0100000011100100: color_data = 12'b001110100111;
		16'b0100000011100101: color_data = 12'b001110100111;
		16'b0100000011100110: color_data = 12'b001110100111;
		16'b0100000011100111: color_data = 12'b001110100111;
		16'b0100000011101000: color_data = 12'b001110100111;
		16'b0100000011101001: color_data = 12'b001110100111;
		16'b0100000011101010: color_data = 12'b001110100111;
		16'b0100000011101011: color_data = 12'b001110100111;
		16'b0100000011101100: color_data = 12'b001110100111;
		16'b0100000011101101: color_data = 12'b001110100111;
		16'b0100000011101110: color_data = 12'b001110100111;
		16'b0100000011101111: color_data = 12'b001110100111;
		16'b0100000011110110: color_data = 12'b001110100111;
		16'b0100000011110111: color_data = 12'b001110100111;
		16'b0100000011111000: color_data = 12'b001110100111;
		16'b0100000011111001: color_data = 12'b001110100111;
		16'b0100000011111010: color_data = 12'b001110100111;
		16'b0100000011111011: color_data = 12'b001110100111;
		16'b0100000011111100: color_data = 12'b001110100111;
		16'b0100000011111101: color_data = 12'b001110100111;
		16'b0100000011111110: color_data = 12'b001110100111;
		16'b0100000011111111: color_data = 12'b001110100111;
		16'b0100000100000000: color_data = 12'b001110100111;
		16'b0100000100000001: color_data = 12'b001110100111;
		16'b0100000100011010: color_data = 12'b001110100111;
		16'b0100000100011011: color_data = 12'b001110100111;
		16'b0100000100011100: color_data = 12'b001110100111;
		16'b0100000100011101: color_data = 12'b001110100111;
		16'b0100000100011110: color_data = 12'b001110100111;
		16'b0100000100011111: color_data = 12'b001110100111;
		16'b0100000100100000: color_data = 12'b001110100111;
		16'b0100000100100001: color_data = 12'b001110100111;
		16'b0100000100100010: color_data = 12'b001110100111;
		16'b0100000100100011: color_data = 12'b001110100111;
		16'b0100000100100100: color_data = 12'b001110100111;
		16'b0100000100100101: color_data = 12'b001110100111;
		16'b0100000100100110: color_data = 12'b001110100111;
		16'b0100000100101101: color_data = 12'b001110100111;
		16'b0100000100101110: color_data = 12'b001110100111;
		16'b0100000100101111: color_data = 12'b001110100111;
		16'b0100000100110000: color_data = 12'b001110100111;
		16'b0100000100110001: color_data = 12'b001110100111;
		16'b0100000100110010: color_data = 12'b001110100111;
		16'b0100000100110011: color_data = 12'b001110100111;
		16'b0100000100110100: color_data = 12'b001110100111;
		16'b0100000100110101: color_data = 12'b001110100111;
		16'b0100000100110110: color_data = 12'b001110100111;
		16'b0100000100110111: color_data = 12'b001110100111;
		16'b0100000100111000: color_data = 12'b001110100111;
		16'b0100000101000101: color_data = 12'b001110100111;
		16'b0100000101000110: color_data = 12'b001110100111;
		16'b0100000101000111: color_data = 12'b001110100111;
		16'b0100000101001000: color_data = 12'b001110100111;
		16'b0100000101001001: color_data = 12'b001110100111;
		16'b0100000101001010: color_data = 12'b001110100111;
		16'b0100000101001011: color_data = 12'b001110100111;
		16'b0100000101001100: color_data = 12'b001110100111;
		16'b0100000101001101: color_data = 12'b001110100111;
		16'b0100000101001110: color_data = 12'b001110100111;
		16'b0100000101001111: color_data = 12'b001110100111;
		16'b0100000101010000: color_data = 12'b001110100111;
		16'b0100000101010001: color_data = 12'b001110100111;
		16'b0100000101011000: color_data = 12'b001110100111;
		16'b0100000101011001: color_data = 12'b001110100111;
		16'b0100000101011010: color_data = 12'b001110100111;
		16'b0100000101011011: color_data = 12'b001110100111;
		16'b0100000101011100: color_data = 12'b001110100111;
		16'b0100000101011101: color_data = 12'b001110100111;
		16'b0100000101011110: color_data = 12'b001110100111;
		16'b0100000101011111: color_data = 12'b001110100111;
		16'b0100000101100000: color_data = 12'b001110100111;
		16'b0100000101100001: color_data = 12'b001110100111;
		16'b0100000101100010: color_data = 12'b001110100111;
		16'b0100000101100011: color_data = 12'b001110100111;
		16'b0100001000000000: color_data = 12'b001110100111;
		16'b0100001000000001: color_data = 12'b001110100111;
		16'b0100001000000010: color_data = 12'b001110100111;
		16'b0100001000000011: color_data = 12'b001110100111;
		16'b0100001000000100: color_data = 12'b001110100111;
		16'b0100001000000101: color_data = 12'b001110100111;
		16'b0100001000000110: color_data = 12'b001110100111;
		16'b0100001000000111: color_data = 12'b001110100111;
		16'b0100001000001000: color_data = 12'b001110100111;
		16'b0100001000001001: color_data = 12'b001110100111;
		16'b0100001000001010: color_data = 12'b001110100111;
		16'b0100001000001011: color_data = 12'b001110100111;
		16'b0100001000001100: color_data = 12'b001110100111;
		16'b0100001000001101: color_data = 12'b001110100111;
		16'b0100001000001110: color_data = 12'b001110100111;
		16'b0100001000001111: color_data = 12'b001110100111;
		16'b0100001000010000: color_data = 12'b001110100111;
		16'b0100001000010001: color_data = 12'b001110100111;
		16'b0100001000010010: color_data = 12'b001110100111;
		16'b0100001000101011: color_data = 12'b001110100111;
		16'b0100001000101100: color_data = 12'b001110100111;
		16'b0100001000101101: color_data = 12'b001110100111;
		16'b0100001000101110: color_data = 12'b001110100111;
		16'b0100001000101111: color_data = 12'b001110100111;
		16'b0100001000110000: color_data = 12'b001110100111;
		16'b0100001000110001: color_data = 12'b001110100111;
		16'b0100001000110010: color_data = 12'b001110100111;
		16'b0100001000110011: color_data = 12'b001110100111;
		16'b0100001000110100: color_data = 12'b001110100111;
		16'b0100001000110101: color_data = 12'b001110100111;
		16'b0100001000110110: color_data = 12'b001110100111;
		16'b0100001000110111: color_data = 12'b001110100111;
		16'b0100001001000100: color_data = 12'b001110100111;
		16'b0100001001000101: color_data = 12'b001110100111;
		16'b0100001001000110: color_data = 12'b001110100111;
		16'b0100001001000111: color_data = 12'b001110100111;
		16'b0100001001001000: color_data = 12'b001110100111;
		16'b0100001001001001: color_data = 12'b001110100111;
		16'b0100001001001010: color_data = 12'b001110100111;
		16'b0100001001001011: color_data = 12'b001110100111;
		16'b0100001001001100: color_data = 12'b001110100111;
		16'b0100001001001101: color_data = 12'b001110100111;
		16'b0100001001001110: color_data = 12'b001110100111;
		16'b0100001001001111: color_data = 12'b001110100111;
		16'b0100001001011100: color_data = 12'b001110100111;
		16'b0100001001011101: color_data = 12'b001110100111;
		16'b0100001001011110: color_data = 12'b001110100111;
		16'b0100001001011111: color_data = 12'b001110100111;
		16'b0100001001100000: color_data = 12'b001110100111;
		16'b0100001001100001: color_data = 12'b001110100111;
		16'b0100001001100010: color_data = 12'b001110100111;
		16'b0100001001100011: color_data = 12'b001110100111;
		16'b0100001001100100: color_data = 12'b001110100111;
		16'b0100001001100101: color_data = 12'b001110100111;
		16'b0100001001100110: color_data = 12'b001110100111;
		16'b0100001001100111: color_data = 12'b001110100111;
		16'b0100001001101000: color_data = 12'b001110100111;
		16'b0100001001110101: color_data = 12'b001110100111;
		16'b0100001001110110: color_data = 12'b001110100111;
		16'b0100001001110111: color_data = 12'b001110100111;
		16'b0100001001111000: color_data = 12'b001110100111;
		16'b0100001001111001: color_data = 12'b001110100111;
		16'b0100001001111010: color_data = 12'b001110100111;
		16'b0100001001111011: color_data = 12'b001110100111;
		16'b0100001001111100: color_data = 12'b001110100111;
		16'b0100001001111101: color_data = 12'b001110100111;
		16'b0100001001111110: color_data = 12'b001110100111;
		16'b0100001001111111: color_data = 12'b001110100111;
		16'b0100001010000000: color_data = 12'b001110100111;
		16'b0100001010001101: color_data = 12'b001110100111;
		16'b0100001010001110: color_data = 12'b001110100111;
		16'b0100001010001111: color_data = 12'b001110100111;
		16'b0100001010010000: color_data = 12'b001110100111;
		16'b0100001010010001: color_data = 12'b001110100111;
		16'b0100001010010010: color_data = 12'b001110100111;
		16'b0100001010010011: color_data = 12'b001110100111;
		16'b0100001010010100: color_data = 12'b001110100111;
		16'b0100001010010101: color_data = 12'b001110100111;
		16'b0100001010010110: color_data = 12'b001110100111;
		16'b0100001010010111: color_data = 12'b001110100111;
		16'b0100001010011000: color_data = 12'b001110100111;
		16'b0100001010011001: color_data = 12'b001110100111;
		16'b0100001010100000: color_data = 12'b001110100111;
		16'b0100001010100001: color_data = 12'b001110100111;
		16'b0100001010100010: color_data = 12'b001110100111;
		16'b0100001010100011: color_data = 12'b001110100111;
		16'b0100001010100100: color_data = 12'b001110100111;
		16'b0100001010100101: color_data = 12'b001110100111;
		16'b0100001010100110: color_data = 12'b001110100111;
		16'b0100001010100111: color_data = 12'b001110100111;
		16'b0100001010101000: color_data = 12'b001110100111;
		16'b0100001010101001: color_data = 12'b001110100111;
		16'b0100001010101010: color_data = 12'b001110100111;
		16'b0100001010101011: color_data = 12'b001110100111;
		16'b0100001011001011: color_data = 12'b001110100111;
		16'b0100001011001100: color_data = 12'b001110100111;
		16'b0100001011001101: color_data = 12'b001110100111;
		16'b0100001011001110: color_data = 12'b001110100111;
		16'b0100001011001111: color_data = 12'b001110100111;
		16'b0100001011010000: color_data = 12'b001110100111;
		16'b0100001011010001: color_data = 12'b001110100111;
		16'b0100001011010010: color_data = 12'b001110100111;
		16'b0100001011010011: color_data = 12'b001110100111;
		16'b0100001011010100: color_data = 12'b001110100111;
		16'b0100001011010101: color_data = 12'b001110100111;
		16'b0100001011010110: color_data = 12'b001110100111;
		16'b0100001011100011: color_data = 12'b001110100111;
		16'b0100001011100100: color_data = 12'b001110100111;
		16'b0100001011100101: color_data = 12'b001110100111;
		16'b0100001011100110: color_data = 12'b001110100111;
		16'b0100001011100111: color_data = 12'b001110100111;
		16'b0100001011101000: color_data = 12'b001110100111;
		16'b0100001011101001: color_data = 12'b001110100111;
		16'b0100001011101010: color_data = 12'b001110100111;
		16'b0100001011101011: color_data = 12'b001110100111;
		16'b0100001011101100: color_data = 12'b001110100111;
		16'b0100001011101101: color_data = 12'b001110100111;
		16'b0100001011101110: color_data = 12'b001110100111;
		16'b0100001011101111: color_data = 12'b001110100111;
		16'b0100001011110110: color_data = 12'b001110100111;
		16'b0100001011110111: color_data = 12'b001110100111;
		16'b0100001011111000: color_data = 12'b001110100111;
		16'b0100001011111001: color_data = 12'b001110100111;
		16'b0100001011111010: color_data = 12'b001110100111;
		16'b0100001011111011: color_data = 12'b001110100111;
		16'b0100001011111100: color_data = 12'b001110100111;
		16'b0100001011111101: color_data = 12'b001110100111;
		16'b0100001011111110: color_data = 12'b001110100111;
		16'b0100001011111111: color_data = 12'b001110100111;
		16'b0100001100000000: color_data = 12'b001110100111;
		16'b0100001100000001: color_data = 12'b001110100111;
		16'b0100001100011010: color_data = 12'b001110100111;
		16'b0100001100011011: color_data = 12'b001110100111;
		16'b0100001100011100: color_data = 12'b001110100111;
		16'b0100001100011101: color_data = 12'b001110100111;
		16'b0100001100011110: color_data = 12'b001110100111;
		16'b0100001100011111: color_data = 12'b001110100111;
		16'b0100001100100000: color_data = 12'b001110100111;
		16'b0100001100100001: color_data = 12'b001110100111;
		16'b0100001100100010: color_data = 12'b001110100111;
		16'b0100001100100011: color_data = 12'b001110100111;
		16'b0100001100100100: color_data = 12'b001110100111;
		16'b0100001100100101: color_data = 12'b001110100111;
		16'b0100001100100110: color_data = 12'b001110100111;
		16'b0100001100101101: color_data = 12'b001110100111;
		16'b0100001100101110: color_data = 12'b001110100111;
		16'b0100001100101111: color_data = 12'b001110100111;
		16'b0100001100110000: color_data = 12'b001110100111;
		16'b0100001100110001: color_data = 12'b001110100111;
		16'b0100001100110010: color_data = 12'b001110100111;
		16'b0100001100110011: color_data = 12'b001110100111;
		16'b0100001100110100: color_data = 12'b001110100111;
		16'b0100001100110101: color_data = 12'b001110100111;
		16'b0100001100110110: color_data = 12'b001110100111;
		16'b0100001100110111: color_data = 12'b001110100111;
		16'b0100001100111000: color_data = 12'b001110100111;
		16'b0100001101000101: color_data = 12'b001110100111;
		16'b0100001101000110: color_data = 12'b001110100111;
		16'b0100001101000111: color_data = 12'b001110100111;
		16'b0100001101001000: color_data = 12'b001110100111;
		16'b0100001101001001: color_data = 12'b001110100111;
		16'b0100001101001010: color_data = 12'b001110100111;
		16'b0100001101001011: color_data = 12'b001110100111;
		16'b0100001101001100: color_data = 12'b001110100111;
		16'b0100001101001101: color_data = 12'b001110100111;
		16'b0100001101001110: color_data = 12'b001110100111;
		16'b0100001101001111: color_data = 12'b001110100111;
		16'b0100001101010000: color_data = 12'b001110100111;
		16'b0100001101010001: color_data = 12'b001110100111;
		16'b0100001101011000: color_data = 12'b001110100111;
		16'b0100001101011001: color_data = 12'b001110100111;
		16'b0100001101011010: color_data = 12'b001110100111;
		16'b0100001101011011: color_data = 12'b001110100111;
		16'b0100001101011100: color_data = 12'b001110100111;
		16'b0100001101011101: color_data = 12'b001110100111;
		16'b0100001101011110: color_data = 12'b001110100111;
		16'b0100001101011111: color_data = 12'b001110100111;
		16'b0100001101100000: color_data = 12'b001110100111;
		16'b0100001101100001: color_data = 12'b001110100111;
		16'b0100001101100010: color_data = 12'b001110100111;
		16'b0100001101100011: color_data = 12'b001110100111;
		16'b0100010000000000: color_data = 12'b001110100111;
		16'b0100010000000001: color_data = 12'b001110100111;
		16'b0100010000000010: color_data = 12'b001110100111;
		16'b0100010000000011: color_data = 12'b001110100111;
		16'b0100010000000100: color_data = 12'b001110100111;
		16'b0100010000000101: color_data = 12'b001110100111;
		16'b0100010000000110: color_data = 12'b001110100111;
		16'b0100010000000111: color_data = 12'b001110100111;
		16'b0100010000001000: color_data = 12'b001110100111;
		16'b0100010000001001: color_data = 12'b001110100111;
		16'b0100010000001010: color_data = 12'b001110100111;
		16'b0100010000001011: color_data = 12'b001110100111;
		16'b0100010000001100: color_data = 12'b001110100111;
		16'b0100010000001101: color_data = 12'b001110100111;
		16'b0100010000001110: color_data = 12'b001110100111;
		16'b0100010000001111: color_data = 12'b001110100111;
		16'b0100010000010000: color_data = 12'b001110100111;
		16'b0100010000010001: color_data = 12'b001110100111;
		16'b0100010000010010: color_data = 12'b001110100111;
		16'b0100010000101011: color_data = 12'b001110100111;
		16'b0100010000101100: color_data = 12'b001110100111;
		16'b0100010000101101: color_data = 12'b001110100111;
		16'b0100010000101110: color_data = 12'b001110100111;
		16'b0100010000101111: color_data = 12'b001110100111;
		16'b0100010000110000: color_data = 12'b001110100111;
		16'b0100010000110001: color_data = 12'b001110100111;
		16'b0100010000110010: color_data = 12'b001110100111;
		16'b0100010000110011: color_data = 12'b001110100111;
		16'b0100010000110100: color_data = 12'b001110100111;
		16'b0100010000110101: color_data = 12'b001110100111;
		16'b0100010000110110: color_data = 12'b001110100111;
		16'b0100010000110111: color_data = 12'b001110100111;
		16'b0100010001000100: color_data = 12'b001110100111;
		16'b0100010001000101: color_data = 12'b001110100111;
		16'b0100010001000110: color_data = 12'b001110100111;
		16'b0100010001000111: color_data = 12'b001110100111;
		16'b0100010001001000: color_data = 12'b001110100111;
		16'b0100010001001001: color_data = 12'b001110100111;
		16'b0100010001001010: color_data = 12'b001110100111;
		16'b0100010001001011: color_data = 12'b001110100111;
		16'b0100010001001100: color_data = 12'b001110100111;
		16'b0100010001001101: color_data = 12'b001110100111;
		16'b0100010001001110: color_data = 12'b001110100111;
		16'b0100010001001111: color_data = 12'b001110100111;
		16'b0100010001011100: color_data = 12'b001110100111;
		16'b0100010001011101: color_data = 12'b001110100111;
		16'b0100010001011110: color_data = 12'b001110100111;
		16'b0100010001011111: color_data = 12'b001110100111;
		16'b0100010001100000: color_data = 12'b001110100111;
		16'b0100010001100001: color_data = 12'b001110100111;
		16'b0100010001100010: color_data = 12'b001110100111;
		16'b0100010001100011: color_data = 12'b001110100111;
		16'b0100010001100100: color_data = 12'b001110100111;
		16'b0100010001100101: color_data = 12'b001110100111;
		16'b0100010001100110: color_data = 12'b001110100111;
		16'b0100010001100111: color_data = 12'b001110100111;
		16'b0100010001101000: color_data = 12'b001110100111;
		16'b0100010001110101: color_data = 12'b001110100111;
		16'b0100010001110110: color_data = 12'b001110100111;
		16'b0100010001110111: color_data = 12'b001110100111;
		16'b0100010001111000: color_data = 12'b001110100111;
		16'b0100010001111001: color_data = 12'b001110100111;
		16'b0100010001111010: color_data = 12'b001110100111;
		16'b0100010001111011: color_data = 12'b001110100111;
		16'b0100010001111100: color_data = 12'b001110100111;
		16'b0100010001111101: color_data = 12'b001110100111;
		16'b0100010001111110: color_data = 12'b001110100111;
		16'b0100010001111111: color_data = 12'b001110100111;
		16'b0100010010000000: color_data = 12'b001110100111;
		16'b0100010010001101: color_data = 12'b001110100111;
		16'b0100010010001110: color_data = 12'b001110100111;
		16'b0100010010001111: color_data = 12'b001110100111;
		16'b0100010010010000: color_data = 12'b001110100111;
		16'b0100010010010001: color_data = 12'b001110100111;
		16'b0100010010010010: color_data = 12'b001110100111;
		16'b0100010010010011: color_data = 12'b001110100111;
		16'b0100010010010100: color_data = 12'b001110100111;
		16'b0100010010010101: color_data = 12'b001110100111;
		16'b0100010010010110: color_data = 12'b001110100111;
		16'b0100010010010111: color_data = 12'b001110100111;
		16'b0100010010011000: color_data = 12'b001110100111;
		16'b0100010010011001: color_data = 12'b001110100111;
		16'b0100010010100000: color_data = 12'b001110100111;
		16'b0100010010100001: color_data = 12'b001110100111;
		16'b0100010010100010: color_data = 12'b001110100111;
		16'b0100010010100011: color_data = 12'b001110100111;
		16'b0100010010100100: color_data = 12'b001110100111;
		16'b0100010010100101: color_data = 12'b001110100111;
		16'b0100010010100110: color_data = 12'b001110100111;
		16'b0100010010100111: color_data = 12'b001110100111;
		16'b0100010010101000: color_data = 12'b001110100111;
		16'b0100010010101001: color_data = 12'b001110100111;
		16'b0100010010101010: color_data = 12'b001110100111;
		16'b0100010010101011: color_data = 12'b001110100111;
		16'b0100010011001011: color_data = 12'b001110100111;
		16'b0100010011001100: color_data = 12'b001110100111;
		16'b0100010011001101: color_data = 12'b001110100111;
		16'b0100010011001110: color_data = 12'b001110100111;
		16'b0100010011001111: color_data = 12'b001110100111;
		16'b0100010011010000: color_data = 12'b001110100111;
		16'b0100010011010001: color_data = 12'b001110100111;
		16'b0100010011010010: color_data = 12'b001110100111;
		16'b0100010011010011: color_data = 12'b001110100111;
		16'b0100010011010100: color_data = 12'b001110100111;
		16'b0100010011010101: color_data = 12'b001110100111;
		16'b0100010011010110: color_data = 12'b001110100111;
		16'b0100010011100011: color_data = 12'b001110100111;
		16'b0100010011100100: color_data = 12'b001110100111;
		16'b0100010011100101: color_data = 12'b001110100111;
		16'b0100010011100110: color_data = 12'b001110100111;
		16'b0100010011100111: color_data = 12'b001110100111;
		16'b0100010011101000: color_data = 12'b001110100111;
		16'b0100010011101001: color_data = 12'b001110100111;
		16'b0100010011101010: color_data = 12'b001110100111;
		16'b0100010011101011: color_data = 12'b001110100111;
		16'b0100010011101100: color_data = 12'b001110100111;
		16'b0100010011101101: color_data = 12'b001110100111;
		16'b0100010011101110: color_data = 12'b001110100111;
		16'b0100010011101111: color_data = 12'b001110100111;
		16'b0100010011110110: color_data = 12'b001110100111;
		16'b0100010011110111: color_data = 12'b001110100111;
		16'b0100010011111000: color_data = 12'b001110100111;
		16'b0100010011111001: color_data = 12'b001110100111;
		16'b0100010011111010: color_data = 12'b001110100111;
		16'b0100010011111011: color_data = 12'b001110100111;
		16'b0100010011111100: color_data = 12'b001110100111;
		16'b0100010011111101: color_data = 12'b001110100111;
		16'b0100010011111110: color_data = 12'b001110100111;
		16'b0100010011111111: color_data = 12'b001110100111;
		16'b0100010100000000: color_data = 12'b001110100111;
		16'b0100010100000001: color_data = 12'b001110100111;
		16'b0100010100011010: color_data = 12'b001110100111;
		16'b0100010100011011: color_data = 12'b001110100111;
		16'b0100010100011100: color_data = 12'b001110100111;
		16'b0100010100011101: color_data = 12'b001110100111;
		16'b0100010100011110: color_data = 12'b001110100111;
		16'b0100010100011111: color_data = 12'b001110100111;
		16'b0100010100100000: color_data = 12'b001110100111;
		16'b0100010100100001: color_data = 12'b001110100111;
		16'b0100010100100010: color_data = 12'b001110100111;
		16'b0100010100100011: color_data = 12'b001110100111;
		16'b0100010100100100: color_data = 12'b001110100111;
		16'b0100010100100101: color_data = 12'b001110100111;
		16'b0100010100100110: color_data = 12'b001110100111;
		16'b0100010100101101: color_data = 12'b001110100111;
		16'b0100010100101110: color_data = 12'b001110100111;
		16'b0100010100101111: color_data = 12'b001110100111;
		16'b0100010100110000: color_data = 12'b001110100111;
		16'b0100010100110001: color_data = 12'b001110100111;
		16'b0100010100110010: color_data = 12'b001110100111;
		16'b0100010100110011: color_data = 12'b001110100111;
		16'b0100010100110100: color_data = 12'b001110100111;
		16'b0100010100110101: color_data = 12'b001110100111;
		16'b0100010100110110: color_data = 12'b001110100111;
		16'b0100010100110111: color_data = 12'b001110100111;
		16'b0100010100111000: color_data = 12'b001110100111;
		16'b0100010101000101: color_data = 12'b001110100111;
		16'b0100010101000110: color_data = 12'b001110100111;
		16'b0100010101000111: color_data = 12'b001110100111;
		16'b0100010101001000: color_data = 12'b001110100111;
		16'b0100010101001001: color_data = 12'b001110100111;
		16'b0100010101001010: color_data = 12'b001110100111;
		16'b0100010101001011: color_data = 12'b001110100111;
		16'b0100010101001100: color_data = 12'b001110100111;
		16'b0100010101001101: color_data = 12'b001110100111;
		16'b0100010101001110: color_data = 12'b001110100111;
		16'b0100010101001111: color_data = 12'b001110100111;
		16'b0100010101010000: color_data = 12'b001110100111;
		16'b0100010101010001: color_data = 12'b001110100111;
		16'b0100010101011000: color_data = 12'b001110100111;
		16'b0100010101011001: color_data = 12'b001110100111;
		16'b0100010101011010: color_data = 12'b001110100111;
		16'b0100010101011011: color_data = 12'b001110100111;
		16'b0100010101011100: color_data = 12'b001110100111;
		16'b0100010101011101: color_data = 12'b001110100111;
		16'b0100010101011110: color_data = 12'b001110100111;
		16'b0100010101011111: color_data = 12'b001110100111;
		16'b0100010101100000: color_data = 12'b001110100111;
		16'b0100010101100001: color_data = 12'b001110100111;
		16'b0100010101100010: color_data = 12'b001110100111;
		16'b0100010101100011: color_data = 12'b001110100111;
		16'b0100011000000000: color_data = 12'b001110100111;
		16'b0100011000000001: color_data = 12'b001110100111;
		16'b0100011000000010: color_data = 12'b001110100111;
		16'b0100011000000011: color_data = 12'b001110100111;
		16'b0100011000000100: color_data = 12'b001110100111;
		16'b0100011000000101: color_data = 12'b001110100111;
		16'b0100011000000110: color_data = 12'b001110100111;
		16'b0100011000000111: color_data = 12'b001110100111;
		16'b0100011000001000: color_data = 12'b001110100111;
		16'b0100011000001001: color_data = 12'b001110100111;
		16'b0100011000001010: color_data = 12'b001110100111;
		16'b0100011000001011: color_data = 12'b001110100111;
		16'b0100011000001100: color_data = 12'b001110100111;
		16'b0100011000001101: color_data = 12'b001110100111;
		16'b0100011000001110: color_data = 12'b001110100111;
		16'b0100011000001111: color_data = 12'b001110100111;
		16'b0100011000010000: color_data = 12'b001110100111;
		16'b0100011000010001: color_data = 12'b001110100111;
		16'b0100011000010010: color_data = 12'b001110100111;
		16'b0100011000101011: color_data = 12'b001110100111;
		16'b0100011000101100: color_data = 12'b001110100111;
		16'b0100011000101101: color_data = 12'b001110100111;
		16'b0100011000101110: color_data = 12'b001110100111;
		16'b0100011000101111: color_data = 12'b001110100111;
		16'b0100011000110000: color_data = 12'b001110100111;
		16'b0100011000110001: color_data = 12'b001110100111;
		16'b0100011000110010: color_data = 12'b001110100111;
		16'b0100011000110011: color_data = 12'b001110100111;
		16'b0100011000110100: color_data = 12'b001110100111;
		16'b0100011000110101: color_data = 12'b001110100111;
		16'b0100011000110110: color_data = 12'b001110100111;
		16'b0100011000110111: color_data = 12'b001110100111;
		16'b0100011001000100: color_data = 12'b001110100111;
		16'b0100011001000101: color_data = 12'b001110100111;
		16'b0100011001000110: color_data = 12'b001110100111;
		16'b0100011001000111: color_data = 12'b001110100111;
		16'b0100011001001000: color_data = 12'b001110100111;
		16'b0100011001001001: color_data = 12'b001110100111;
		16'b0100011001001010: color_data = 12'b001110100111;
		16'b0100011001001011: color_data = 12'b001110100111;
		16'b0100011001001100: color_data = 12'b001110100111;
		16'b0100011001001101: color_data = 12'b001110100111;
		16'b0100011001001110: color_data = 12'b001110100111;
		16'b0100011001001111: color_data = 12'b001110100111;
		16'b0100011001011100: color_data = 12'b001110100111;
		16'b0100011001011101: color_data = 12'b001110100111;
		16'b0100011001011110: color_data = 12'b001110100111;
		16'b0100011001011111: color_data = 12'b001110100111;
		16'b0100011001100000: color_data = 12'b001110100111;
		16'b0100011001100001: color_data = 12'b001110100111;
		16'b0100011001100010: color_data = 12'b001110100111;
		16'b0100011001100011: color_data = 12'b001110100111;
		16'b0100011001100100: color_data = 12'b001110100111;
		16'b0100011001100101: color_data = 12'b001110100111;
		16'b0100011001100110: color_data = 12'b001110100111;
		16'b0100011001100111: color_data = 12'b001110100111;
		16'b0100011001101000: color_data = 12'b001110100111;
		16'b0100011001110101: color_data = 12'b001110100111;
		16'b0100011001110110: color_data = 12'b001110100111;
		16'b0100011001110111: color_data = 12'b001110100111;
		16'b0100011001111000: color_data = 12'b001110100111;
		16'b0100011001111001: color_data = 12'b001110100111;
		16'b0100011001111010: color_data = 12'b001110100111;
		16'b0100011001111011: color_data = 12'b001110100111;
		16'b0100011001111100: color_data = 12'b001110100111;
		16'b0100011001111101: color_data = 12'b001110100111;
		16'b0100011001111110: color_data = 12'b001110100111;
		16'b0100011001111111: color_data = 12'b001110100111;
		16'b0100011010000000: color_data = 12'b001110100111;
		16'b0100011010001101: color_data = 12'b001110100111;
		16'b0100011010001110: color_data = 12'b001110100111;
		16'b0100011010001111: color_data = 12'b001110100111;
		16'b0100011010010000: color_data = 12'b001110100111;
		16'b0100011010010001: color_data = 12'b001110100111;
		16'b0100011010010010: color_data = 12'b001110100111;
		16'b0100011010010011: color_data = 12'b001110100111;
		16'b0100011010010100: color_data = 12'b001110100111;
		16'b0100011010010101: color_data = 12'b001110100111;
		16'b0100011010010110: color_data = 12'b001110100111;
		16'b0100011010010111: color_data = 12'b001110100111;
		16'b0100011010011000: color_data = 12'b001110100111;
		16'b0100011010011001: color_data = 12'b001110100111;
		16'b0100011010100000: color_data = 12'b001110100111;
		16'b0100011010100001: color_data = 12'b001110100111;
		16'b0100011010100010: color_data = 12'b001110100111;
		16'b0100011010100011: color_data = 12'b001110100111;
		16'b0100011010100100: color_data = 12'b001110100111;
		16'b0100011010100101: color_data = 12'b001110100111;
		16'b0100011010100110: color_data = 12'b001110100111;
		16'b0100011010100111: color_data = 12'b001110100111;
		16'b0100011010101000: color_data = 12'b001110100111;
		16'b0100011010101001: color_data = 12'b001110100111;
		16'b0100011010101010: color_data = 12'b001110100111;
		16'b0100011010101011: color_data = 12'b001110100111;
		16'b0100011011001011: color_data = 12'b001110100111;
		16'b0100011011001100: color_data = 12'b001110100111;
		16'b0100011011001101: color_data = 12'b001110100111;
		16'b0100011011001110: color_data = 12'b001110100111;
		16'b0100011011001111: color_data = 12'b001110100111;
		16'b0100011011010000: color_data = 12'b001110100111;
		16'b0100011011010001: color_data = 12'b001110100111;
		16'b0100011011010010: color_data = 12'b001110100111;
		16'b0100011011010011: color_data = 12'b001110100111;
		16'b0100011011010100: color_data = 12'b001110100111;
		16'b0100011011010101: color_data = 12'b001110100111;
		16'b0100011011010110: color_data = 12'b001110100111;
		16'b0100011011100011: color_data = 12'b001110100111;
		16'b0100011011100100: color_data = 12'b001110100111;
		16'b0100011011100101: color_data = 12'b001110100111;
		16'b0100011011100110: color_data = 12'b001110100111;
		16'b0100011011100111: color_data = 12'b001110100111;
		16'b0100011011101000: color_data = 12'b001110100111;
		16'b0100011011101001: color_data = 12'b001110100111;
		16'b0100011011101010: color_data = 12'b001110100111;
		16'b0100011011101011: color_data = 12'b001110100111;
		16'b0100011011101100: color_data = 12'b001110100111;
		16'b0100011011101101: color_data = 12'b001110100111;
		16'b0100011011101110: color_data = 12'b001110100111;
		16'b0100011011101111: color_data = 12'b001110100111;
		16'b0100011011110110: color_data = 12'b001110100111;
		16'b0100011011110111: color_data = 12'b001110100111;
		16'b0100011011111000: color_data = 12'b001110100111;
		16'b0100011011111001: color_data = 12'b001110100111;
		16'b0100011011111010: color_data = 12'b001110100111;
		16'b0100011011111011: color_data = 12'b001110100111;
		16'b0100011011111100: color_data = 12'b001110100111;
		16'b0100011011111101: color_data = 12'b001110100111;
		16'b0100011011111110: color_data = 12'b001110100111;
		16'b0100011011111111: color_data = 12'b001110100111;
		16'b0100011100000000: color_data = 12'b001110100111;
		16'b0100011100000001: color_data = 12'b001110100111;
		16'b0100011100011010: color_data = 12'b001110100111;
		16'b0100011100011011: color_data = 12'b001110100111;
		16'b0100011100011100: color_data = 12'b001110100111;
		16'b0100011100011101: color_data = 12'b001110100111;
		16'b0100011100011110: color_data = 12'b001110100111;
		16'b0100011100011111: color_data = 12'b001110100111;
		16'b0100011100100000: color_data = 12'b001110100111;
		16'b0100011100100001: color_data = 12'b001110100111;
		16'b0100011100100010: color_data = 12'b001110100111;
		16'b0100011100100011: color_data = 12'b001110100111;
		16'b0100011100100100: color_data = 12'b001110100111;
		16'b0100011100100101: color_data = 12'b001110100111;
		16'b0100011100100110: color_data = 12'b001110100111;
		16'b0100011100101101: color_data = 12'b001110100111;
		16'b0100011100101110: color_data = 12'b001110100111;
		16'b0100011100101111: color_data = 12'b001110100111;
		16'b0100011100110000: color_data = 12'b001110100111;
		16'b0100011100110001: color_data = 12'b001110100111;
		16'b0100011100110010: color_data = 12'b001110100111;
		16'b0100011100110011: color_data = 12'b001110100111;
		16'b0100011100110100: color_data = 12'b001110100111;
		16'b0100011100110101: color_data = 12'b001110100111;
		16'b0100011100110110: color_data = 12'b001110100111;
		16'b0100011100110111: color_data = 12'b001110100111;
		16'b0100011100111000: color_data = 12'b001110100111;
		16'b0100011101000101: color_data = 12'b001110100111;
		16'b0100011101000110: color_data = 12'b001110100111;
		16'b0100011101000111: color_data = 12'b001110100111;
		16'b0100011101001000: color_data = 12'b001110100111;
		16'b0100011101001001: color_data = 12'b001110100111;
		16'b0100011101001010: color_data = 12'b001110100111;
		16'b0100011101001011: color_data = 12'b001110100111;
		16'b0100011101001100: color_data = 12'b001110100111;
		16'b0100011101001101: color_data = 12'b001110100111;
		16'b0100011101001110: color_data = 12'b001110100111;
		16'b0100011101001111: color_data = 12'b001110100111;
		16'b0100011101010000: color_data = 12'b001110100111;
		16'b0100011101010001: color_data = 12'b001110100111;
		16'b0100011101011000: color_data = 12'b001110100111;
		16'b0100011101011001: color_data = 12'b001110100111;
		16'b0100011101011010: color_data = 12'b001110100111;
		16'b0100011101011011: color_data = 12'b001110100111;
		16'b0100011101011100: color_data = 12'b001110100111;
		16'b0100011101011101: color_data = 12'b001110100111;
		16'b0100011101011110: color_data = 12'b001110100111;
		16'b0100011101011111: color_data = 12'b001110100111;
		16'b0100011101100000: color_data = 12'b001110100111;
		16'b0100011101100001: color_data = 12'b001110100111;
		16'b0100011101100010: color_data = 12'b001110100111;
		16'b0100011101100011: color_data = 12'b001110100111;
		16'b0100100000000000: color_data = 12'b001110100111;
		16'b0100100000000001: color_data = 12'b001110100111;
		16'b0100100000000010: color_data = 12'b001110100111;
		16'b0100100000000011: color_data = 12'b001110100111;
		16'b0100100000000100: color_data = 12'b001110100111;
		16'b0100100000000101: color_data = 12'b001110100111;
		16'b0100100000000110: color_data = 12'b001110100111;
		16'b0100100000000111: color_data = 12'b001110100111;
		16'b0100100000001000: color_data = 12'b001110100111;
		16'b0100100000001001: color_data = 12'b001110100111;
		16'b0100100000001010: color_data = 12'b001110100111;
		16'b0100100000001011: color_data = 12'b001110100111;
		16'b0100100000001100: color_data = 12'b001110100111;
		16'b0100100000001101: color_data = 12'b001110100111;
		16'b0100100000001110: color_data = 12'b001110100111;
		16'b0100100000001111: color_data = 12'b001110100111;
		16'b0100100000010000: color_data = 12'b001110100111;
		16'b0100100000010001: color_data = 12'b001110100111;
		16'b0100100000010010: color_data = 12'b001110100111;
		16'b0100100000101011: color_data = 12'b001110100111;
		16'b0100100000101100: color_data = 12'b001110100111;
		16'b0100100000101101: color_data = 12'b001110100111;
		16'b0100100000101110: color_data = 12'b001110100111;
		16'b0100100000101111: color_data = 12'b001110100111;
		16'b0100100000110000: color_data = 12'b001110100111;
		16'b0100100000110001: color_data = 12'b001110100111;
		16'b0100100000110010: color_data = 12'b001110100111;
		16'b0100100000110011: color_data = 12'b001110100111;
		16'b0100100000110100: color_data = 12'b001110100111;
		16'b0100100000110101: color_data = 12'b001110100111;
		16'b0100100000110110: color_data = 12'b001110100111;
		16'b0100100000110111: color_data = 12'b001110100111;
		16'b0100100001000100: color_data = 12'b001110100111;
		16'b0100100001000101: color_data = 12'b001110100111;
		16'b0100100001000110: color_data = 12'b001110100111;
		16'b0100100001000111: color_data = 12'b001110100111;
		16'b0100100001001000: color_data = 12'b001110100111;
		16'b0100100001001001: color_data = 12'b001110100111;
		16'b0100100001001010: color_data = 12'b001110100111;
		16'b0100100001001011: color_data = 12'b001110100111;
		16'b0100100001001100: color_data = 12'b001110100111;
		16'b0100100001001101: color_data = 12'b001110100111;
		16'b0100100001001110: color_data = 12'b001110100111;
		16'b0100100001001111: color_data = 12'b001110100111;
		16'b0100100001011100: color_data = 12'b001110100111;
		16'b0100100001011101: color_data = 12'b001110100111;
		16'b0100100001011110: color_data = 12'b001110100111;
		16'b0100100001011111: color_data = 12'b001110100111;
		16'b0100100001100000: color_data = 12'b001110100111;
		16'b0100100001100001: color_data = 12'b001110100111;
		16'b0100100001100010: color_data = 12'b001110100111;
		16'b0100100001100011: color_data = 12'b001110100111;
		16'b0100100001100100: color_data = 12'b001110100111;
		16'b0100100001100101: color_data = 12'b001110100111;
		16'b0100100001100110: color_data = 12'b001110100111;
		16'b0100100001100111: color_data = 12'b001110100111;
		16'b0100100001101000: color_data = 12'b001110100111;
		16'b0100100001110101: color_data = 12'b001110100111;
		16'b0100100001110110: color_data = 12'b001110100111;
		16'b0100100001110111: color_data = 12'b001110100111;
		16'b0100100001111000: color_data = 12'b001110100111;
		16'b0100100001111001: color_data = 12'b001110100111;
		16'b0100100001111010: color_data = 12'b001110100111;
		16'b0100100001111011: color_data = 12'b001110100111;
		16'b0100100001111100: color_data = 12'b001110100111;
		16'b0100100001111101: color_data = 12'b001110100111;
		16'b0100100001111110: color_data = 12'b001110100111;
		16'b0100100001111111: color_data = 12'b001110100111;
		16'b0100100010000000: color_data = 12'b001110100111;
		16'b0100100010001101: color_data = 12'b001110100111;
		16'b0100100010001110: color_data = 12'b001110100111;
		16'b0100100010001111: color_data = 12'b001110100111;
		16'b0100100010010000: color_data = 12'b001110100111;
		16'b0100100010010001: color_data = 12'b001110100111;
		16'b0100100010010010: color_data = 12'b001110100111;
		16'b0100100010010011: color_data = 12'b001110100111;
		16'b0100100010010100: color_data = 12'b001110100111;
		16'b0100100010010101: color_data = 12'b001110100111;
		16'b0100100010010110: color_data = 12'b001110100111;
		16'b0100100010010111: color_data = 12'b001110100111;
		16'b0100100010011000: color_data = 12'b001110100111;
		16'b0100100010011001: color_data = 12'b001110100111;
		16'b0100100010100000: color_data = 12'b001110100111;
		16'b0100100010100001: color_data = 12'b001110100111;
		16'b0100100010100010: color_data = 12'b001110100111;
		16'b0100100010100011: color_data = 12'b001110100111;
		16'b0100100010100100: color_data = 12'b001110100111;
		16'b0100100010100101: color_data = 12'b001110100111;
		16'b0100100010100110: color_data = 12'b001110100111;
		16'b0100100010100111: color_data = 12'b001110100111;
		16'b0100100010101000: color_data = 12'b001110100111;
		16'b0100100010101001: color_data = 12'b001110100111;
		16'b0100100010101010: color_data = 12'b001110100111;
		16'b0100100010101011: color_data = 12'b001110100111;
		16'b0100100011001011: color_data = 12'b001110100111;
		16'b0100100011001100: color_data = 12'b001110100111;
		16'b0100100011001101: color_data = 12'b001110100111;
		16'b0100100011001110: color_data = 12'b001110100111;
		16'b0100100011001111: color_data = 12'b001110100111;
		16'b0100100011010000: color_data = 12'b001110100111;
		16'b0100100011010001: color_data = 12'b001110100111;
		16'b0100100011010010: color_data = 12'b001110100111;
		16'b0100100011010011: color_data = 12'b001110100111;
		16'b0100100011010100: color_data = 12'b001110100111;
		16'b0100100011010101: color_data = 12'b001110100111;
		16'b0100100011010110: color_data = 12'b001110100111;
		16'b0100100011100011: color_data = 12'b001110100111;
		16'b0100100011100100: color_data = 12'b001110100111;
		16'b0100100011100101: color_data = 12'b001110100111;
		16'b0100100011100110: color_data = 12'b001110100111;
		16'b0100100011100111: color_data = 12'b001110100111;
		16'b0100100011101000: color_data = 12'b001110100111;
		16'b0100100011101001: color_data = 12'b001110100111;
		16'b0100100011101010: color_data = 12'b001110100111;
		16'b0100100011101011: color_data = 12'b001110100111;
		16'b0100100011101100: color_data = 12'b001110100111;
		16'b0100100011101101: color_data = 12'b001110100111;
		16'b0100100011101110: color_data = 12'b001110100111;
		16'b0100100011101111: color_data = 12'b001110100111;
		16'b0100100011110110: color_data = 12'b001110100111;
		16'b0100100011110111: color_data = 12'b001110100111;
		16'b0100100011111000: color_data = 12'b001110100111;
		16'b0100100011111001: color_data = 12'b001110100111;
		16'b0100100011111010: color_data = 12'b001110100111;
		16'b0100100011111011: color_data = 12'b001110100111;
		16'b0100100011111100: color_data = 12'b001110100111;
		16'b0100100011111101: color_data = 12'b001110100111;
		16'b0100100011111110: color_data = 12'b001110100111;
		16'b0100100011111111: color_data = 12'b001110100111;
		16'b0100100100000000: color_data = 12'b001110100111;
		16'b0100100100000001: color_data = 12'b001110100111;
		16'b0100100100011010: color_data = 12'b001110100111;
		16'b0100100100011011: color_data = 12'b001110100111;
		16'b0100100100011100: color_data = 12'b001110100111;
		16'b0100100100011101: color_data = 12'b001110100111;
		16'b0100100100011110: color_data = 12'b001110100111;
		16'b0100100100011111: color_data = 12'b001110100111;
		16'b0100100100100000: color_data = 12'b001110100111;
		16'b0100100100100001: color_data = 12'b001110100111;
		16'b0100100100100010: color_data = 12'b001110100111;
		16'b0100100100100011: color_data = 12'b001110100111;
		16'b0100100100100100: color_data = 12'b001110100111;
		16'b0100100100100101: color_data = 12'b001110100111;
		16'b0100100100100110: color_data = 12'b001110100111;
		16'b0100100100101101: color_data = 12'b001110100111;
		16'b0100100100101110: color_data = 12'b001110100111;
		16'b0100100100101111: color_data = 12'b001110100111;
		16'b0100100100110000: color_data = 12'b001110100111;
		16'b0100100100110001: color_data = 12'b001110100111;
		16'b0100100100110010: color_data = 12'b001110100111;
		16'b0100100100110011: color_data = 12'b001110100111;
		16'b0100100100110100: color_data = 12'b001110100111;
		16'b0100100100110101: color_data = 12'b001110100111;
		16'b0100100100110110: color_data = 12'b001110100111;
		16'b0100100100110111: color_data = 12'b001110100111;
		16'b0100100100111000: color_data = 12'b001110100111;
		16'b0100100101000101: color_data = 12'b001110100111;
		16'b0100100101000110: color_data = 12'b001110100111;
		16'b0100100101000111: color_data = 12'b001110100111;
		16'b0100100101001000: color_data = 12'b001110100111;
		16'b0100100101001001: color_data = 12'b001110100111;
		16'b0100100101001010: color_data = 12'b001110100111;
		16'b0100100101001011: color_data = 12'b001110100111;
		16'b0100100101001100: color_data = 12'b001110100111;
		16'b0100100101001101: color_data = 12'b001110100111;
		16'b0100100101001110: color_data = 12'b001110100111;
		16'b0100100101001111: color_data = 12'b001110100111;
		16'b0100100101010000: color_data = 12'b001110100111;
		16'b0100100101010001: color_data = 12'b001110100111;
		16'b0100100101011000: color_data = 12'b001110100111;
		16'b0100100101011001: color_data = 12'b001110100111;
		16'b0100100101011010: color_data = 12'b001110100111;
		16'b0100100101011011: color_data = 12'b001110100111;
		16'b0100100101011100: color_data = 12'b001110100111;
		16'b0100100101011101: color_data = 12'b001110100111;
		16'b0100100101011110: color_data = 12'b001110100111;
		16'b0100100101011111: color_data = 12'b001110100111;
		16'b0100100101100000: color_data = 12'b001110100111;
		16'b0100100101100001: color_data = 12'b001110100111;
		16'b0100100101100010: color_data = 12'b001110100111;
		16'b0100100101100011: color_data = 12'b001110100111;
		16'b0100101000000000: color_data = 12'b001110100111;
		16'b0100101000000001: color_data = 12'b001110100111;
		16'b0100101000000010: color_data = 12'b001110100111;
		16'b0100101000000011: color_data = 12'b001110100111;
		16'b0100101000000100: color_data = 12'b001110100111;
		16'b0100101000000101: color_data = 12'b001110100111;
		16'b0100101000000110: color_data = 12'b001110100111;
		16'b0100101000000111: color_data = 12'b001110100111;
		16'b0100101000001000: color_data = 12'b001110100111;
		16'b0100101000001001: color_data = 12'b001110100111;
		16'b0100101000001010: color_data = 12'b001110100111;
		16'b0100101000001011: color_data = 12'b001110100111;
		16'b0100101000001100: color_data = 12'b001110100111;
		16'b0100101000001101: color_data = 12'b001110100111;
		16'b0100101000001110: color_data = 12'b001110100111;
		16'b0100101000001111: color_data = 12'b001110100111;
		16'b0100101000010000: color_data = 12'b001110100111;
		16'b0100101000010001: color_data = 12'b001110100111;
		16'b0100101000010010: color_data = 12'b001110100111;
		16'b0100101000101011: color_data = 12'b001110100111;
		16'b0100101000101100: color_data = 12'b001110100111;
		16'b0100101000101101: color_data = 12'b001110100111;
		16'b0100101000101110: color_data = 12'b001110100111;
		16'b0100101000101111: color_data = 12'b001110100111;
		16'b0100101000110000: color_data = 12'b001110100111;
		16'b0100101000110001: color_data = 12'b001110100111;
		16'b0100101000110010: color_data = 12'b001110100111;
		16'b0100101000110011: color_data = 12'b001110100111;
		16'b0100101000110100: color_data = 12'b001110100111;
		16'b0100101000110101: color_data = 12'b001110100111;
		16'b0100101000110110: color_data = 12'b001110100111;
		16'b0100101000110111: color_data = 12'b001110100111;
		16'b0100101001000100: color_data = 12'b001110100111;
		16'b0100101001000101: color_data = 12'b001110100111;
		16'b0100101001000110: color_data = 12'b001110100111;
		16'b0100101001000111: color_data = 12'b001110100111;
		16'b0100101001001000: color_data = 12'b001110100111;
		16'b0100101001001001: color_data = 12'b001110100111;
		16'b0100101001001010: color_data = 12'b001110100111;
		16'b0100101001001011: color_data = 12'b001110100111;
		16'b0100101001001100: color_data = 12'b001110100111;
		16'b0100101001001101: color_data = 12'b001110100111;
		16'b0100101001001110: color_data = 12'b001110100111;
		16'b0100101001001111: color_data = 12'b001110100111;
		16'b0100101001011100: color_data = 12'b001110100111;
		16'b0100101001011101: color_data = 12'b001110100111;
		16'b0100101001011110: color_data = 12'b001110100111;
		16'b0100101001011111: color_data = 12'b001110100111;
		16'b0100101001100000: color_data = 12'b001110100111;
		16'b0100101001100001: color_data = 12'b001110100111;
		16'b0100101001100010: color_data = 12'b001110100111;
		16'b0100101001100011: color_data = 12'b001110100111;
		16'b0100101001100100: color_data = 12'b001110100111;
		16'b0100101001100101: color_data = 12'b001110100111;
		16'b0100101001100110: color_data = 12'b001110100111;
		16'b0100101001100111: color_data = 12'b001110100111;
		16'b0100101001101000: color_data = 12'b001110100111;
		16'b0100101001110101: color_data = 12'b001110100111;
		16'b0100101001110110: color_data = 12'b001110100111;
		16'b0100101001110111: color_data = 12'b001110100111;
		16'b0100101001111000: color_data = 12'b001110100111;
		16'b0100101001111001: color_data = 12'b001110100111;
		16'b0100101001111010: color_data = 12'b001110100111;
		16'b0100101001111011: color_data = 12'b001110100111;
		16'b0100101001111100: color_data = 12'b001110100111;
		16'b0100101001111101: color_data = 12'b001110100111;
		16'b0100101001111110: color_data = 12'b001110100111;
		16'b0100101001111111: color_data = 12'b001110100111;
		16'b0100101010000000: color_data = 12'b001110100111;
		16'b0100101010001101: color_data = 12'b001110100111;
		16'b0100101010001110: color_data = 12'b001110100111;
		16'b0100101010001111: color_data = 12'b001110100111;
		16'b0100101010010000: color_data = 12'b001110100111;
		16'b0100101010010001: color_data = 12'b001110100111;
		16'b0100101010010010: color_data = 12'b001110100111;
		16'b0100101010010011: color_data = 12'b001110100111;
		16'b0100101010010100: color_data = 12'b001110100111;
		16'b0100101010010101: color_data = 12'b001110100111;
		16'b0100101010010110: color_data = 12'b001110100111;
		16'b0100101010010111: color_data = 12'b001110100111;
		16'b0100101010011000: color_data = 12'b001110100111;
		16'b0100101010011001: color_data = 12'b001110100111;
		16'b0100101010100000: color_data = 12'b001110100111;
		16'b0100101010100001: color_data = 12'b001110100111;
		16'b0100101010100010: color_data = 12'b001110100111;
		16'b0100101010100011: color_data = 12'b001110100111;
		16'b0100101010100100: color_data = 12'b001110100111;
		16'b0100101010100101: color_data = 12'b001110100111;
		16'b0100101010100110: color_data = 12'b001110100111;
		16'b0100101010100111: color_data = 12'b001110100111;
		16'b0100101010101000: color_data = 12'b001110100111;
		16'b0100101010101001: color_data = 12'b001110100111;
		16'b0100101010101010: color_data = 12'b001110100111;
		16'b0100101010101011: color_data = 12'b001110100111;
		16'b0100101011001011: color_data = 12'b001110100111;
		16'b0100101011001100: color_data = 12'b001110100111;
		16'b0100101011001101: color_data = 12'b001110100111;
		16'b0100101011001110: color_data = 12'b001110100111;
		16'b0100101011001111: color_data = 12'b001110100111;
		16'b0100101011010000: color_data = 12'b001110100111;
		16'b0100101011010001: color_data = 12'b001110100111;
		16'b0100101011010010: color_data = 12'b001110100111;
		16'b0100101011010011: color_data = 12'b001110100111;
		16'b0100101011010100: color_data = 12'b001110100111;
		16'b0100101011010101: color_data = 12'b001110100111;
		16'b0100101011010110: color_data = 12'b001110100111;
		16'b0100101011100011: color_data = 12'b001110100111;
		16'b0100101011100100: color_data = 12'b001110100111;
		16'b0100101011100101: color_data = 12'b001110100111;
		16'b0100101011100110: color_data = 12'b001110100111;
		16'b0100101011100111: color_data = 12'b001110100111;
		16'b0100101011101000: color_data = 12'b001110100111;
		16'b0100101011101001: color_data = 12'b001110100111;
		16'b0100101011101010: color_data = 12'b001110100111;
		16'b0100101011101011: color_data = 12'b001110100111;
		16'b0100101011101100: color_data = 12'b001110100111;
		16'b0100101011101101: color_data = 12'b001110100111;
		16'b0100101011101110: color_data = 12'b001110100111;
		16'b0100101011101111: color_data = 12'b001110100111;
		16'b0100101011110110: color_data = 12'b001110100111;
		16'b0100101011110111: color_data = 12'b001110100111;
		16'b0100101011111000: color_data = 12'b001110100111;
		16'b0100101011111001: color_data = 12'b001110100111;
		16'b0100101011111010: color_data = 12'b001110100111;
		16'b0100101011111011: color_data = 12'b001110100111;
		16'b0100101011111100: color_data = 12'b001110100111;
		16'b0100101011111101: color_data = 12'b001110100111;
		16'b0100101011111110: color_data = 12'b001110100111;
		16'b0100101011111111: color_data = 12'b001110100111;
		16'b0100101100000000: color_data = 12'b001110100111;
		16'b0100101100000001: color_data = 12'b001110100111;
		16'b0100101100011010: color_data = 12'b001110100111;
		16'b0100101100011011: color_data = 12'b001110100111;
		16'b0100101100011100: color_data = 12'b001110100111;
		16'b0100101100011101: color_data = 12'b001110100111;
		16'b0100101100011110: color_data = 12'b001110100111;
		16'b0100101100011111: color_data = 12'b001110100111;
		16'b0100101100100000: color_data = 12'b001110100111;
		16'b0100101100100001: color_data = 12'b001110100111;
		16'b0100101100100010: color_data = 12'b001110100111;
		16'b0100101100100011: color_data = 12'b001110100111;
		16'b0100101100100100: color_data = 12'b001110100111;
		16'b0100101100100101: color_data = 12'b001110100111;
		16'b0100101100100110: color_data = 12'b001110100111;
		16'b0100101100101101: color_data = 12'b001110100111;
		16'b0100101100101110: color_data = 12'b001110100111;
		16'b0100101100101111: color_data = 12'b001110100111;
		16'b0100101100110000: color_data = 12'b001110100111;
		16'b0100101100110001: color_data = 12'b001110100111;
		16'b0100101100110010: color_data = 12'b001110100111;
		16'b0100101100110011: color_data = 12'b001110100111;
		16'b0100101100110100: color_data = 12'b001110100111;
		16'b0100101100110101: color_data = 12'b001110100111;
		16'b0100101100110110: color_data = 12'b001110100111;
		16'b0100101100110111: color_data = 12'b001110100111;
		16'b0100101100111000: color_data = 12'b001110100111;
		16'b0100101101000101: color_data = 12'b001110100111;
		16'b0100101101000110: color_data = 12'b001110100111;
		16'b0100101101000111: color_data = 12'b001110100111;
		16'b0100101101001000: color_data = 12'b001110100111;
		16'b0100101101001001: color_data = 12'b001110100111;
		16'b0100101101001010: color_data = 12'b001110100111;
		16'b0100101101001011: color_data = 12'b001110100111;
		16'b0100101101001100: color_data = 12'b001110100111;
		16'b0100101101001101: color_data = 12'b001110100111;
		16'b0100101101001110: color_data = 12'b001110100111;
		16'b0100101101001111: color_data = 12'b001110100111;
		16'b0100101101010000: color_data = 12'b001110100111;
		16'b0100101101010001: color_data = 12'b001110100111;
		16'b0100101101011000: color_data = 12'b001110100111;
		16'b0100101101011001: color_data = 12'b001110100111;
		16'b0100101101011010: color_data = 12'b001110100111;
		16'b0100101101011011: color_data = 12'b001110100111;
		16'b0100101101011100: color_data = 12'b001110100111;
		16'b0100101101011101: color_data = 12'b001110100111;
		16'b0100101101011110: color_data = 12'b001110100111;
		16'b0100101101011111: color_data = 12'b001110100111;
		16'b0100101101100000: color_data = 12'b001110100111;
		16'b0100101101100001: color_data = 12'b001110100111;
		16'b0100101101100010: color_data = 12'b001110100111;
		16'b0100101101100011: color_data = 12'b001110100111;
		16'b0100110000000000: color_data = 12'b001110100111;
		16'b0100110000000001: color_data = 12'b001110100111;
		16'b0100110000000010: color_data = 12'b001110100111;
		16'b0100110000000011: color_data = 12'b001110100111;
		16'b0100110000000100: color_data = 12'b001110100111;
		16'b0100110000000101: color_data = 12'b001110100111;
		16'b0100110000000110: color_data = 12'b001110100111;
		16'b0100110000000111: color_data = 12'b001110100111;
		16'b0100110000001000: color_data = 12'b001110100111;
		16'b0100110000001001: color_data = 12'b001110100111;
		16'b0100110000001010: color_data = 12'b001110100111;
		16'b0100110000001011: color_data = 12'b001110100111;
		16'b0100110000001100: color_data = 12'b001110100111;
		16'b0100110000101011: color_data = 12'b001110100111;
		16'b0100110000101100: color_data = 12'b001110100111;
		16'b0100110000101101: color_data = 12'b001110100111;
		16'b0100110000101110: color_data = 12'b001110100111;
		16'b0100110000101111: color_data = 12'b001110100111;
		16'b0100110000110000: color_data = 12'b001110100111;
		16'b0100110000110001: color_data = 12'b001110100111;
		16'b0100110000110010: color_data = 12'b001110100111;
		16'b0100110000110011: color_data = 12'b001110100111;
		16'b0100110000110100: color_data = 12'b001110100111;
		16'b0100110000110101: color_data = 12'b001110100111;
		16'b0100110000110110: color_data = 12'b001110100111;
		16'b0100110000110111: color_data = 12'b001110100111;
		16'b0100110000111000: color_data = 12'b001110100111;
		16'b0100110000111001: color_data = 12'b001110100111;
		16'b0100110000111010: color_data = 12'b001110100111;
		16'b0100110000111011: color_data = 12'b001110100111;
		16'b0100110000111100: color_data = 12'b001110100111;
		16'b0100110000111101: color_data = 12'b001110100111;
		16'b0100110000111110: color_data = 12'b001110100111;
		16'b0100110000111111: color_data = 12'b001110100111;
		16'b0100110001000000: color_data = 12'b001110100111;
		16'b0100110001000001: color_data = 12'b001110100111;
		16'b0100110001000010: color_data = 12'b001110100111;
		16'b0100110001000011: color_data = 12'b001110100111;
		16'b0100110001000100: color_data = 12'b001110100111;
		16'b0100110001000101: color_data = 12'b001110100111;
		16'b0100110001000110: color_data = 12'b001110100111;
		16'b0100110001000111: color_data = 12'b001110100111;
		16'b0100110001001000: color_data = 12'b001110100111;
		16'b0100110001001001: color_data = 12'b001110100111;
		16'b0100110001001010: color_data = 12'b001110100111;
		16'b0100110001001011: color_data = 12'b001110100111;
		16'b0100110001001100: color_data = 12'b001110100111;
		16'b0100110001001101: color_data = 12'b001110100111;
		16'b0100110001001110: color_data = 12'b001110100111;
		16'b0100110001001111: color_data = 12'b001110100111;
		16'b0100110001011100: color_data = 12'b001110100111;
		16'b0100110001011101: color_data = 12'b001110100111;
		16'b0100110001011110: color_data = 12'b001110100111;
		16'b0100110001011111: color_data = 12'b001110100111;
		16'b0100110001100000: color_data = 12'b001110100111;
		16'b0100110001100001: color_data = 12'b001110100111;
		16'b0100110001100010: color_data = 12'b001110100111;
		16'b0100110001100011: color_data = 12'b001110100111;
		16'b0100110001100100: color_data = 12'b001110100111;
		16'b0100110001100101: color_data = 12'b001110100111;
		16'b0100110001100110: color_data = 12'b001110100111;
		16'b0100110001100111: color_data = 12'b001110100111;
		16'b0100110001101000: color_data = 12'b001110100111;
		16'b0100110001110101: color_data = 12'b001110100111;
		16'b0100110001110110: color_data = 12'b001110100111;
		16'b0100110001110111: color_data = 12'b001110100111;
		16'b0100110001111000: color_data = 12'b001110100111;
		16'b0100110001111001: color_data = 12'b001110100111;
		16'b0100110001111010: color_data = 12'b001110100111;
		16'b0100110001111011: color_data = 12'b001110100111;
		16'b0100110001111100: color_data = 12'b001110100111;
		16'b0100110001111101: color_data = 12'b001110100111;
		16'b0100110001111110: color_data = 12'b001110100111;
		16'b0100110001111111: color_data = 12'b001110100111;
		16'b0100110010000000: color_data = 12'b001110100111;
		16'b0100110010001101: color_data = 12'b001110100111;
		16'b0100110010001110: color_data = 12'b001110100111;
		16'b0100110010001111: color_data = 12'b001110100111;
		16'b0100110010010000: color_data = 12'b001110100111;
		16'b0100110010010001: color_data = 12'b001110100111;
		16'b0100110010010010: color_data = 12'b001110100111;
		16'b0100110010010011: color_data = 12'b001110100111;
		16'b0100110010010100: color_data = 12'b001110100111;
		16'b0100110010010101: color_data = 12'b001110100111;
		16'b0100110010010110: color_data = 12'b001110100111;
		16'b0100110010010111: color_data = 12'b001110100111;
		16'b0100110010011000: color_data = 12'b001110100111;
		16'b0100110010011001: color_data = 12'b001110100111;
		16'b0100110010100000: color_data = 12'b001110100111;
		16'b0100110010100001: color_data = 12'b001110100111;
		16'b0100110010100010: color_data = 12'b001110100111;
		16'b0100110010100011: color_data = 12'b001110100111;
		16'b0100110010100100: color_data = 12'b001110100111;
		16'b0100110010100101: color_data = 12'b001110100111;
		16'b0100110010100110: color_data = 12'b001110100111;
		16'b0100110010100111: color_data = 12'b001110100111;
		16'b0100110010101000: color_data = 12'b001110100111;
		16'b0100110010101001: color_data = 12'b001110100111;
		16'b0100110010101010: color_data = 12'b001110100111;
		16'b0100110010101011: color_data = 12'b001110100111;
		16'b0100110011001011: color_data = 12'b001110100111;
		16'b0100110011001100: color_data = 12'b001110100111;
		16'b0100110011001101: color_data = 12'b001110100111;
		16'b0100110011001110: color_data = 12'b001110100111;
		16'b0100110011001111: color_data = 12'b001110100111;
		16'b0100110011010000: color_data = 12'b001110100111;
		16'b0100110011010001: color_data = 12'b001110100111;
		16'b0100110011010010: color_data = 12'b001110100111;
		16'b0100110011010011: color_data = 12'b001110100111;
		16'b0100110011010100: color_data = 12'b001110100111;
		16'b0100110011010101: color_data = 12'b001110100111;
		16'b0100110011010110: color_data = 12'b001110100111;
		16'b0100110011010111: color_data = 12'b001110100111;
		16'b0100110011011000: color_data = 12'b001110100111;
		16'b0100110011011001: color_data = 12'b001110100111;
		16'b0100110011011010: color_data = 12'b001110100111;
		16'b0100110011011011: color_data = 12'b001110100111;
		16'b0100110011011100: color_data = 12'b001110100111;
		16'b0100110011011101: color_data = 12'b001110100111;
		16'b0100110011011110: color_data = 12'b001110100111;
		16'b0100110011011111: color_data = 12'b001110100111;
		16'b0100110011100000: color_data = 12'b001110100111;
		16'b0100110011100001: color_data = 12'b001110100111;
		16'b0100110011100010: color_data = 12'b001110100111;
		16'b0100110011100011: color_data = 12'b001110100111;
		16'b0100110011100100: color_data = 12'b001110100111;
		16'b0100110011100101: color_data = 12'b001110100111;
		16'b0100110011100110: color_data = 12'b001110100111;
		16'b0100110011100111: color_data = 12'b001110100111;
		16'b0100110011101000: color_data = 12'b001110100111;
		16'b0100110011110110: color_data = 12'b001110100111;
		16'b0100110011110111: color_data = 12'b001110100111;
		16'b0100110011111000: color_data = 12'b001110100111;
		16'b0100110011111001: color_data = 12'b001110100111;
		16'b0100110011111010: color_data = 12'b001110100111;
		16'b0100110011111011: color_data = 12'b001110100111;
		16'b0100110011111100: color_data = 12'b001110100111;
		16'b0100110011111101: color_data = 12'b001110100111;
		16'b0100110011111110: color_data = 12'b001110100111;
		16'b0100110011111111: color_data = 12'b001110100111;
		16'b0100110100000000: color_data = 12'b001110100111;
		16'b0100110100000001: color_data = 12'b001110100111;
		16'b0100110100011010: color_data = 12'b001110100111;
		16'b0100110100011011: color_data = 12'b001110100111;
		16'b0100110100011100: color_data = 12'b001110100111;
		16'b0100110100011101: color_data = 12'b001110100111;
		16'b0100110100011110: color_data = 12'b001110100111;
		16'b0100110100011111: color_data = 12'b001110100111;
		16'b0100110100100000: color_data = 12'b001110100111;
		16'b0100110100100001: color_data = 12'b001110100111;
		16'b0100110100100010: color_data = 12'b001110100111;
		16'b0100110100100011: color_data = 12'b001110100111;
		16'b0100110100100100: color_data = 12'b001110100111;
		16'b0100110100100101: color_data = 12'b001110100111;
		16'b0100110100100110: color_data = 12'b001110100111;
		16'b0100110100101101: color_data = 12'b001110100111;
		16'b0100110100101110: color_data = 12'b001110100111;
		16'b0100110100101111: color_data = 12'b001110100111;
		16'b0100110100110000: color_data = 12'b001110100111;
		16'b0100110100110001: color_data = 12'b001110100111;
		16'b0100110100110010: color_data = 12'b001110100111;
		16'b0100110100110011: color_data = 12'b001110100111;
		16'b0100110100110100: color_data = 12'b001110100111;
		16'b0100110100110101: color_data = 12'b001110100111;
		16'b0100110100110110: color_data = 12'b001110100111;
		16'b0100110100110111: color_data = 12'b001110100111;
		16'b0100110100111000: color_data = 12'b001110100111;
		16'b0100110101000101: color_data = 12'b001110100111;
		16'b0100110101000110: color_data = 12'b001110100111;
		16'b0100110101000111: color_data = 12'b001110100111;
		16'b0100110101001000: color_data = 12'b001110100111;
		16'b0100110101001001: color_data = 12'b001110100111;
		16'b0100110101001010: color_data = 12'b001110100111;
		16'b0100110101001011: color_data = 12'b001110100111;
		16'b0100110101001100: color_data = 12'b001110100111;
		16'b0100110101001101: color_data = 12'b001110100111;
		16'b0100110101001110: color_data = 12'b001110100111;
		16'b0100110101001111: color_data = 12'b001110100111;
		16'b0100110101010000: color_data = 12'b001110100111;
		16'b0100110101010001: color_data = 12'b001110100111;
		16'b0100110101011000: color_data = 12'b001110100111;
		16'b0100110101011001: color_data = 12'b001110100111;
		16'b0100110101011010: color_data = 12'b001110100111;
		16'b0100110101011011: color_data = 12'b001110100111;
		16'b0100110101011100: color_data = 12'b001110100111;
		16'b0100110101011101: color_data = 12'b001110100111;
		16'b0100110101011110: color_data = 12'b001110100111;
		16'b0100110101011111: color_data = 12'b001110100111;
		16'b0100110101100000: color_data = 12'b001110100111;
		16'b0100110101100001: color_data = 12'b001110100111;
		16'b0100110101100010: color_data = 12'b001110100111;
		16'b0100110101100011: color_data = 12'b001110100111;
		16'b0100111000000000: color_data = 12'b001110100111;
		16'b0100111000000001: color_data = 12'b001110100111;
		16'b0100111000000010: color_data = 12'b001110100111;
		16'b0100111000000011: color_data = 12'b001110100111;
		16'b0100111000000100: color_data = 12'b001110100111;
		16'b0100111000000101: color_data = 12'b001110100111;
		16'b0100111000000110: color_data = 12'b001110100111;
		16'b0100111000000111: color_data = 12'b001110100111;
		16'b0100111000001000: color_data = 12'b001110100111;
		16'b0100111000001001: color_data = 12'b001110100111;
		16'b0100111000001010: color_data = 12'b001110100111;
		16'b0100111000001011: color_data = 12'b001110100111;
		16'b0100111000001100: color_data = 12'b001110100111;
		16'b0100111000101011: color_data = 12'b001110100111;
		16'b0100111000101100: color_data = 12'b001110100111;
		16'b0100111000101101: color_data = 12'b001110100111;
		16'b0100111000101110: color_data = 12'b001110100111;
		16'b0100111000101111: color_data = 12'b001110100111;
		16'b0100111000110000: color_data = 12'b001110100111;
		16'b0100111000110001: color_data = 12'b001110100111;
		16'b0100111000110010: color_data = 12'b001110100111;
		16'b0100111000110011: color_data = 12'b001110100111;
		16'b0100111000110100: color_data = 12'b001110100111;
		16'b0100111000110101: color_data = 12'b001110100111;
		16'b0100111000110110: color_data = 12'b001110100111;
		16'b0100111000110111: color_data = 12'b001110100111;
		16'b0100111000111000: color_data = 12'b001110100111;
		16'b0100111000111001: color_data = 12'b001110100111;
		16'b0100111000111010: color_data = 12'b001110100111;
		16'b0100111000111011: color_data = 12'b001110100111;
		16'b0100111000111100: color_data = 12'b001110100111;
		16'b0100111000111101: color_data = 12'b001110100111;
		16'b0100111000111110: color_data = 12'b001110100111;
		16'b0100111000111111: color_data = 12'b001110100111;
		16'b0100111001000000: color_data = 12'b001110100111;
		16'b0100111001000001: color_data = 12'b001110100111;
		16'b0100111001000010: color_data = 12'b001110100111;
		16'b0100111001000011: color_data = 12'b001110100111;
		16'b0100111001000100: color_data = 12'b001110100111;
		16'b0100111001000101: color_data = 12'b001110100111;
		16'b0100111001000110: color_data = 12'b001110100111;
		16'b0100111001000111: color_data = 12'b001110100111;
		16'b0100111001001000: color_data = 12'b001110100111;
		16'b0100111001001001: color_data = 12'b001110100111;
		16'b0100111001001010: color_data = 12'b001110100111;
		16'b0100111001001011: color_data = 12'b001110100111;
		16'b0100111001001100: color_data = 12'b001110100111;
		16'b0100111001001101: color_data = 12'b001110100111;
		16'b0100111001001110: color_data = 12'b001110100111;
		16'b0100111001001111: color_data = 12'b001110100111;
		16'b0100111001011100: color_data = 12'b001110100111;
		16'b0100111001011101: color_data = 12'b001110100111;
		16'b0100111001011110: color_data = 12'b001110100111;
		16'b0100111001011111: color_data = 12'b001110100111;
		16'b0100111001100000: color_data = 12'b001110100111;
		16'b0100111001100001: color_data = 12'b001110100111;
		16'b0100111001100010: color_data = 12'b001110100111;
		16'b0100111001100011: color_data = 12'b001110100111;
		16'b0100111001100100: color_data = 12'b001110100111;
		16'b0100111001100101: color_data = 12'b001110100111;
		16'b0100111001100110: color_data = 12'b001110100111;
		16'b0100111001100111: color_data = 12'b001110100111;
		16'b0100111001101000: color_data = 12'b001110100111;
		16'b0100111001110101: color_data = 12'b001110100111;
		16'b0100111001110110: color_data = 12'b001110100111;
		16'b0100111001110111: color_data = 12'b001110100111;
		16'b0100111001111000: color_data = 12'b001110100111;
		16'b0100111001111001: color_data = 12'b001110100111;
		16'b0100111001111010: color_data = 12'b001110100111;
		16'b0100111001111011: color_data = 12'b001110100111;
		16'b0100111001111100: color_data = 12'b001110100111;
		16'b0100111001111101: color_data = 12'b001110100111;
		16'b0100111001111110: color_data = 12'b001110100111;
		16'b0100111001111111: color_data = 12'b001110100111;
		16'b0100111010000000: color_data = 12'b001110100111;
		16'b0100111010001101: color_data = 12'b001110100111;
		16'b0100111010001110: color_data = 12'b001110100111;
		16'b0100111010001111: color_data = 12'b001110100111;
		16'b0100111010010000: color_data = 12'b001110100111;
		16'b0100111010010001: color_data = 12'b001110100111;
		16'b0100111010010010: color_data = 12'b001110100111;
		16'b0100111010010011: color_data = 12'b001110100111;
		16'b0100111010010100: color_data = 12'b001110100111;
		16'b0100111010010101: color_data = 12'b001110100111;
		16'b0100111010010110: color_data = 12'b001110100111;
		16'b0100111010010111: color_data = 12'b001110100111;
		16'b0100111010011000: color_data = 12'b001110100111;
		16'b0100111010011001: color_data = 12'b001110100111;
		16'b0100111010100000: color_data = 12'b001110100111;
		16'b0100111010100001: color_data = 12'b001110100111;
		16'b0100111010100010: color_data = 12'b001110100111;
		16'b0100111010100011: color_data = 12'b001110100111;
		16'b0100111010100100: color_data = 12'b001110100111;
		16'b0100111010100101: color_data = 12'b001110100111;
		16'b0100111010100110: color_data = 12'b001110100111;
		16'b0100111010100111: color_data = 12'b001110100111;
		16'b0100111010101000: color_data = 12'b001110100111;
		16'b0100111010101001: color_data = 12'b001110100111;
		16'b0100111010101010: color_data = 12'b001110100111;
		16'b0100111010101011: color_data = 12'b001110100111;
		16'b0100111011001011: color_data = 12'b001110100111;
		16'b0100111011001100: color_data = 12'b001110100111;
		16'b0100111011001101: color_data = 12'b001110100111;
		16'b0100111011001110: color_data = 12'b001110100111;
		16'b0100111011001111: color_data = 12'b001110100111;
		16'b0100111011010000: color_data = 12'b001110100111;
		16'b0100111011010001: color_data = 12'b001110100111;
		16'b0100111011010010: color_data = 12'b001110100111;
		16'b0100111011010011: color_data = 12'b001110100111;
		16'b0100111011010100: color_data = 12'b001110100111;
		16'b0100111011010101: color_data = 12'b001110100111;
		16'b0100111011010110: color_data = 12'b001110100111;
		16'b0100111011010111: color_data = 12'b001110100111;
		16'b0100111011011000: color_data = 12'b001110100111;
		16'b0100111011011001: color_data = 12'b001110100111;
		16'b0100111011011010: color_data = 12'b001110100111;
		16'b0100111011011011: color_data = 12'b001110100111;
		16'b0100111011011100: color_data = 12'b001110100111;
		16'b0100111011011101: color_data = 12'b001110100111;
		16'b0100111011011110: color_data = 12'b001110100111;
		16'b0100111011011111: color_data = 12'b001110100111;
		16'b0100111011100000: color_data = 12'b001110100111;
		16'b0100111011100001: color_data = 12'b001110100111;
		16'b0100111011100010: color_data = 12'b001110100111;
		16'b0100111011100011: color_data = 12'b001110100111;
		16'b0100111011100100: color_data = 12'b001110100111;
		16'b0100111011100101: color_data = 12'b001110100111;
		16'b0100111011100110: color_data = 12'b001110100111;
		16'b0100111011100111: color_data = 12'b001110100111;
		16'b0100111011101000: color_data = 12'b001110100111;
		16'b0100111011110110: color_data = 12'b001110100111;
		16'b0100111011110111: color_data = 12'b001110100111;
		16'b0100111011111000: color_data = 12'b001110100111;
		16'b0100111011111001: color_data = 12'b001110100111;
		16'b0100111011111010: color_data = 12'b001110100111;
		16'b0100111011111011: color_data = 12'b001110100111;
		16'b0100111011111100: color_data = 12'b001110100111;
		16'b0100111011111101: color_data = 12'b001110100111;
		16'b0100111011111110: color_data = 12'b001110100111;
		16'b0100111011111111: color_data = 12'b001110100111;
		16'b0100111100000000: color_data = 12'b001110100111;
		16'b0100111100000001: color_data = 12'b001110100111;
		16'b0100111100011010: color_data = 12'b001110100111;
		16'b0100111100011011: color_data = 12'b001110100111;
		16'b0100111100011100: color_data = 12'b001110100111;
		16'b0100111100011101: color_data = 12'b001110100111;
		16'b0100111100011110: color_data = 12'b001110100111;
		16'b0100111100011111: color_data = 12'b001110100111;
		16'b0100111100100000: color_data = 12'b001110100111;
		16'b0100111100100001: color_data = 12'b001110100111;
		16'b0100111100100010: color_data = 12'b001110100111;
		16'b0100111100100011: color_data = 12'b001110100111;
		16'b0100111100100100: color_data = 12'b001110100111;
		16'b0100111100100101: color_data = 12'b001110100111;
		16'b0100111100100110: color_data = 12'b001110100111;
		16'b0100111100101101: color_data = 12'b001110100111;
		16'b0100111100101110: color_data = 12'b001110100111;
		16'b0100111100101111: color_data = 12'b001110100111;
		16'b0100111100110000: color_data = 12'b001110100111;
		16'b0100111100110001: color_data = 12'b001110100111;
		16'b0100111100110010: color_data = 12'b001110100111;
		16'b0100111100110011: color_data = 12'b001110100111;
		16'b0100111100110100: color_data = 12'b001110100111;
		16'b0100111100110101: color_data = 12'b001110100111;
		16'b0100111100110110: color_data = 12'b001110100111;
		16'b0100111100110111: color_data = 12'b001110100111;
		16'b0100111100111000: color_data = 12'b001110100111;
		16'b0100111101000101: color_data = 12'b001110100111;
		16'b0100111101000110: color_data = 12'b001110100111;
		16'b0100111101000111: color_data = 12'b001110100111;
		16'b0100111101001000: color_data = 12'b001110100111;
		16'b0100111101001001: color_data = 12'b001110100111;
		16'b0100111101001010: color_data = 12'b001110100111;
		16'b0100111101001011: color_data = 12'b001110100111;
		16'b0100111101001100: color_data = 12'b001110100111;
		16'b0100111101001101: color_data = 12'b001110100111;
		16'b0100111101001110: color_data = 12'b001110100111;
		16'b0100111101001111: color_data = 12'b001110100111;
		16'b0100111101010000: color_data = 12'b001110100111;
		16'b0100111101010001: color_data = 12'b001110100111;
		16'b0100111101011000: color_data = 12'b001110100111;
		16'b0100111101011001: color_data = 12'b001110100111;
		16'b0100111101011010: color_data = 12'b001110100111;
		16'b0100111101011011: color_data = 12'b001110100111;
		16'b0100111101011100: color_data = 12'b001110100111;
		16'b0100111101011101: color_data = 12'b001110100111;
		16'b0100111101011110: color_data = 12'b001110100111;
		16'b0100111101011111: color_data = 12'b001110100111;
		16'b0100111101100000: color_data = 12'b001110100111;
		16'b0100111101100001: color_data = 12'b001110100111;
		16'b0100111101100010: color_data = 12'b001110100111;
		16'b0100111101100011: color_data = 12'b001110100111;
		16'b0101000000000000: color_data = 12'b001110100111;
		16'b0101000000000001: color_data = 12'b001110100111;
		16'b0101000000000010: color_data = 12'b001110100111;
		16'b0101000000000011: color_data = 12'b001110100111;
		16'b0101000000000100: color_data = 12'b001110100111;
		16'b0101000000000101: color_data = 12'b001110100111;
		16'b0101000000000110: color_data = 12'b001110100111;
		16'b0101000000000111: color_data = 12'b001110100111;
		16'b0101000000001000: color_data = 12'b001110100111;
		16'b0101000000001001: color_data = 12'b001110100111;
		16'b0101000000001010: color_data = 12'b001110100111;
		16'b0101000000001011: color_data = 12'b001110100111;
		16'b0101000000001100: color_data = 12'b001110100111;
		16'b0101000000101011: color_data = 12'b001110100111;
		16'b0101000000101100: color_data = 12'b001110100111;
		16'b0101000000101101: color_data = 12'b001110100111;
		16'b0101000000101110: color_data = 12'b001110100111;
		16'b0101000000101111: color_data = 12'b001110100111;
		16'b0101000000110000: color_data = 12'b001110100111;
		16'b0101000000110001: color_data = 12'b001110100111;
		16'b0101000000110010: color_data = 12'b001110100111;
		16'b0101000000110011: color_data = 12'b001110100111;
		16'b0101000000110100: color_data = 12'b001110100111;
		16'b0101000000110101: color_data = 12'b001110100111;
		16'b0101000000110110: color_data = 12'b001110100111;
		16'b0101000000110111: color_data = 12'b001110100111;
		16'b0101000000111000: color_data = 12'b001110100111;
		16'b0101000000111001: color_data = 12'b001110100111;
		16'b0101000000111010: color_data = 12'b001110100111;
		16'b0101000000111011: color_data = 12'b001110100111;
		16'b0101000000111100: color_data = 12'b001110100111;
		16'b0101000000111101: color_data = 12'b001110100111;
		16'b0101000000111110: color_data = 12'b001110100111;
		16'b0101000000111111: color_data = 12'b001110100111;
		16'b0101000001000000: color_data = 12'b001110100111;
		16'b0101000001000001: color_data = 12'b001110100111;
		16'b0101000001000010: color_data = 12'b001110100111;
		16'b0101000001000011: color_data = 12'b001110100111;
		16'b0101000001000100: color_data = 12'b001110100111;
		16'b0101000001000101: color_data = 12'b001110100111;
		16'b0101000001000110: color_data = 12'b001110100111;
		16'b0101000001000111: color_data = 12'b001110100111;
		16'b0101000001001000: color_data = 12'b001110100111;
		16'b0101000001001001: color_data = 12'b001110100111;
		16'b0101000001001010: color_data = 12'b001110100111;
		16'b0101000001001011: color_data = 12'b001110100111;
		16'b0101000001001100: color_data = 12'b001110100111;
		16'b0101000001001101: color_data = 12'b001110100111;
		16'b0101000001001110: color_data = 12'b001110100111;
		16'b0101000001001111: color_data = 12'b001110100111;
		16'b0101000001011100: color_data = 12'b001110100111;
		16'b0101000001011101: color_data = 12'b001110100111;
		16'b0101000001011110: color_data = 12'b001110100111;
		16'b0101000001011111: color_data = 12'b001110100111;
		16'b0101000001100000: color_data = 12'b001110100111;
		16'b0101000001100001: color_data = 12'b001110100111;
		16'b0101000001100010: color_data = 12'b001110100111;
		16'b0101000001100011: color_data = 12'b001110100111;
		16'b0101000001100100: color_data = 12'b001110100111;
		16'b0101000001100101: color_data = 12'b001110100111;
		16'b0101000001100110: color_data = 12'b001110100111;
		16'b0101000001100111: color_data = 12'b001110100111;
		16'b0101000001101000: color_data = 12'b001110100111;
		16'b0101000001110101: color_data = 12'b001110100111;
		16'b0101000001110110: color_data = 12'b001110100111;
		16'b0101000001110111: color_data = 12'b001110100111;
		16'b0101000001111000: color_data = 12'b001110100111;
		16'b0101000001111001: color_data = 12'b001110100111;
		16'b0101000001111010: color_data = 12'b001110100111;
		16'b0101000001111011: color_data = 12'b001110100111;
		16'b0101000001111100: color_data = 12'b001110100111;
		16'b0101000001111101: color_data = 12'b001110100111;
		16'b0101000001111110: color_data = 12'b001110100111;
		16'b0101000001111111: color_data = 12'b001110100111;
		16'b0101000010000000: color_data = 12'b001110100111;
		16'b0101000010001101: color_data = 12'b001110100111;
		16'b0101000010001110: color_data = 12'b001110100111;
		16'b0101000010001111: color_data = 12'b001110100111;
		16'b0101000010010000: color_data = 12'b001110100111;
		16'b0101000010010001: color_data = 12'b001110100111;
		16'b0101000010010010: color_data = 12'b001110100111;
		16'b0101000010010011: color_data = 12'b001110100111;
		16'b0101000010010100: color_data = 12'b001110100111;
		16'b0101000010010101: color_data = 12'b001110100111;
		16'b0101000010010110: color_data = 12'b001110100111;
		16'b0101000010010111: color_data = 12'b001110100111;
		16'b0101000010011000: color_data = 12'b001110100111;
		16'b0101000010011001: color_data = 12'b001110100111;
		16'b0101000010100000: color_data = 12'b001110100111;
		16'b0101000010100001: color_data = 12'b001110100111;
		16'b0101000010100010: color_data = 12'b001110100111;
		16'b0101000010100011: color_data = 12'b001110100111;
		16'b0101000010100100: color_data = 12'b001110100111;
		16'b0101000010100101: color_data = 12'b001110100111;
		16'b0101000010100110: color_data = 12'b001110100111;
		16'b0101000010100111: color_data = 12'b001110100111;
		16'b0101000010101000: color_data = 12'b001110100111;
		16'b0101000010101001: color_data = 12'b001110100111;
		16'b0101000010101010: color_data = 12'b001110100111;
		16'b0101000010101011: color_data = 12'b001110100111;
		16'b0101000011001011: color_data = 12'b001110100111;
		16'b0101000011001100: color_data = 12'b001110100111;
		16'b0101000011001101: color_data = 12'b001110100111;
		16'b0101000011001110: color_data = 12'b001110100111;
		16'b0101000011001111: color_data = 12'b001110100111;
		16'b0101000011010000: color_data = 12'b001110100111;
		16'b0101000011010001: color_data = 12'b001110100111;
		16'b0101000011010010: color_data = 12'b001110100111;
		16'b0101000011010011: color_data = 12'b001110100111;
		16'b0101000011010100: color_data = 12'b001110100111;
		16'b0101000011010101: color_data = 12'b001110100111;
		16'b0101000011010110: color_data = 12'b001110100111;
		16'b0101000011010111: color_data = 12'b001110100111;
		16'b0101000011011000: color_data = 12'b001110100111;
		16'b0101000011011001: color_data = 12'b001110100111;
		16'b0101000011011010: color_data = 12'b001110100111;
		16'b0101000011011011: color_data = 12'b001110100111;
		16'b0101000011011100: color_data = 12'b001110100111;
		16'b0101000011011101: color_data = 12'b001110100111;
		16'b0101000011011110: color_data = 12'b001110100111;
		16'b0101000011011111: color_data = 12'b001110100111;
		16'b0101000011100000: color_data = 12'b001110100111;
		16'b0101000011100001: color_data = 12'b001110100111;
		16'b0101000011100010: color_data = 12'b001110100111;
		16'b0101000011100011: color_data = 12'b001110100111;
		16'b0101000011100100: color_data = 12'b001110100111;
		16'b0101000011100101: color_data = 12'b001110100111;
		16'b0101000011100110: color_data = 12'b001110100111;
		16'b0101000011100111: color_data = 12'b001110100111;
		16'b0101000011101000: color_data = 12'b001110100111;
		16'b0101000011110110: color_data = 12'b001110100111;
		16'b0101000011110111: color_data = 12'b001110100111;
		16'b0101000011111000: color_data = 12'b001110100111;
		16'b0101000011111001: color_data = 12'b001110100111;
		16'b0101000011111010: color_data = 12'b001110100111;
		16'b0101000011111011: color_data = 12'b001110100111;
		16'b0101000011111100: color_data = 12'b001110100111;
		16'b0101000011111101: color_data = 12'b001110100111;
		16'b0101000011111110: color_data = 12'b001110100111;
		16'b0101000011111111: color_data = 12'b001110100111;
		16'b0101000100000000: color_data = 12'b001110100111;
		16'b0101000100000001: color_data = 12'b001110100111;
		16'b0101000100011010: color_data = 12'b001110100111;
		16'b0101000100011011: color_data = 12'b001110100111;
		16'b0101000100011100: color_data = 12'b001110100111;
		16'b0101000100011101: color_data = 12'b001110100111;
		16'b0101000100011110: color_data = 12'b001110100111;
		16'b0101000100011111: color_data = 12'b001110100111;
		16'b0101000100100000: color_data = 12'b001110100111;
		16'b0101000100100001: color_data = 12'b001110100111;
		16'b0101000100100010: color_data = 12'b001110100111;
		16'b0101000100100011: color_data = 12'b001110100111;
		16'b0101000100100100: color_data = 12'b001110100111;
		16'b0101000100100101: color_data = 12'b001110100111;
		16'b0101000100100110: color_data = 12'b001110100111;
		16'b0101000100101101: color_data = 12'b001110100111;
		16'b0101000100101110: color_data = 12'b001110100111;
		16'b0101000100101111: color_data = 12'b001110100111;
		16'b0101000100110000: color_data = 12'b001110100111;
		16'b0101000100110001: color_data = 12'b001110100111;
		16'b0101000100110010: color_data = 12'b001110100111;
		16'b0101000100110011: color_data = 12'b001110100111;
		16'b0101000100110100: color_data = 12'b001110100111;
		16'b0101000100110101: color_data = 12'b001110100111;
		16'b0101000100110110: color_data = 12'b001110100111;
		16'b0101000100110111: color_data = 12'b001110100111;
		16'b0101000100111000: color_data = 12'b001110100111;
		16'b0101000101000101: color_data = 12'b001110100111;
		16'b0101000101000110: color_data = 12'b001110100111;
		16'b0101000101000111: color_data = 12'b001110100111;
		16'b0101000101001000: color_data = 12'b001110100111;
		16'b0101000101001001: color_data = 12'b001110100111;
		16'b0101000101001010: color_data = 12'b001110100111;
		16'b0101000101001011: color_data = 12'b001110100111;
		16'b0101000101001100: color_data = 12'b001110100111;
		16'b0101000101001101: color_data = 12'b001110100111;
		16'b0101000101001110: color_data = 12'b001110100111;
		16'b0101000101001111: color_data = 12'b001110100111;
		16'b0101000101010000: color_data = 12'b001110100111;
		16'b0101000101010001: color_data = 12'b001110100111;
		16'b0101000101011000: color_data = 12'b001110100111;
		16'b0101000101011001: color_data = 12'b001110100111;
		16'b0101000101011010: color_data = 12'b001110100111;
		16'b0101000101011011: color_data = 12'b001110100111;
		16'b0101000101011100: color_data = 12'b001110100111;
		16'b0101000101011101: color_data = 12'b001110100111;
		16'b0101000101011110: color_data = 12'b001110100111;
		16'b0101000101011111: color_data = 12'b001110100111;
		16'b0101000101100000: color_data = 12'b001110100111;
		16'b0101000101100001: color_data = 12'b001110100111;
		16'b0101000101100010: color_data = 12'b001110100111;
		16'b0101000101100011: color_data = 12'b001110100111;
		16'b0101001000000000: color_data = 12'b001110100111;
		16'b0101001000000001: color_data = 12'b001110100111;
		16'b0101001000000010: color_data = 12'b001110100111;
		16'b0101001000000011: color_data = 12'b001110100111;
		16'b0101001000000100: color_data = 12'b001110100111;
		16'b0101001000000101: color_data = 12'b001110100111;
		16'b0101001000000110: color_data = 12'b001110100111;
		16'b0101001000000111: color_data = 12'b001110100111;
		16'b0101001000001000: color_data = 12'b001110100111;
		16'b0101001000001001: color_data = 12'b001110100111;
		16'b0101001000001010: color_data = 12'b001110100111;
		16'b0101001000001011: color_data = 12'b001110100111;
		16'b0101001000001100: color_data = 12'b001110100111;
		16'b0101001000101011: color_data = 12'b001110100111;
		16'b0101001000101100: color_data = 12'b001110100111;
		16'b0101001000101101: color_data = 12'b001110100111;
		16'b0101001000101110: color_data = 12'b001110100111;
		16'b0101001000101111: color_data = 12'b001110100111;
		16'b0101001000110000: color_data = 12'b001110100111;
		16'b0101001000110001: color_data = 12'b001110100111;
		16'b0101001000110010: color_data = 12'b001110100111;
		16'b0101001000110011: color_data = 12'b001110100111;
		16'b0101001000110100: color_data = 12'b001110100111;
		16'b0101001000110101: color_data = 12'b001110100111;
		16'b0101001000110110: color_data = 12'b001110100111;
		16'b0101001000110111: color_data = 12'b001110100111;
		16'b0101001000111000: color_data = 12'b001110100111;
		16'b0101001000111001: color_data = 12'b001110100111;
		16'b0101001000111010: color_data = 12'b001110100111;
		16'b0101001000111011: color_data = 12'b001110100111;
		16'b0101001000111100: color_data = 12'b001110100111;
		16'b0101001000111101: color_data = 12'b001110100111;
		16'b0101001000111110: color_data = 12'b001110100111;
		16'b0101001000111111: color_data = 12'b001110100111;
		16'b0101001001000000: color_data = 12'b001110100111;
		16'b0101001001000001: color_data = 12'b001110100111;
		16'b0101001001000010: color_data = 12'b001110100111;
		16'b0101001001000011: color_data = 12'b001110100111;
		16'b0101001001000100: color_data = 12'b001110100111;
		16'b0101001001000101: color_data = 12'b001110100111;
		16'b0101001001000110: color_data = 12'b001110100111;
		16'b0101001001000111: color_data = 12'b001110100111;
		16'b0101001001001000: color_data = 12'b001110100111;
		16'b0101001001001001: color_data = 12'b001110100111;
		16'b0101001001001010: color_data = 12'b001110100111;
		16'b0101001001001011: color_data = 12'b001110100111;
		16'b0101001001001100: color_data = 12'b001110100111;
		16'b0101001001001101: color_data = 12'b001110100111;
		16'b0101001001001110: color_data = 12'b001110100111;
		16'b0101001001001111: color_data = 12'b001110100111;
		16'b0101001001011100: color_data = 12'b001110100111;
		16'b0101001001011101: color_data = 12'b001110100111;
		16'b0101001001011110: color_data = 12'b001110100111;
		16'b0101001001011111: color_data = 12'b001110100111;
		16'b0101001001100000: color_data = 12'b001110100111;
		16'b0101001001100001: color_data = 12'b001110100111;
		16'b0101001001100010: color_data = 12'b001110100111;
		16'b0101001001100011: color_data = 12'b001110100111;
		16'b0101001001100100: color_data = 12'b001110100111;
		16'b0101001001100101: color_data = 12'b001110100111;
		16'b0101001001100110: color_data = 12'b001110100111;
		16'b0101001001100111: color_data = 12'b001110100111;
		16'b0101001001101000: color_data = 12'b001110100111;
		16'b0101001001110101: color_data = 12'b001110100111;
		16'b0101001001110110: color_data = 12'b001110100111;
		16'b0101001001110111: color_data = 12'b001110100111;
		16'b0101001001111000: color_data = 12'b001110100111;
		16'b0101001001111001: color_data = 12'b001110100111;
		16'b0101001001111010: color_data = 12'b001110100111;
		16'b0101001001111011: color_data = 12'b001110100111;
		16'b0101001001111100: color_data = 12'b001110100111;
		16'b0101001001111101: color_data = 12'b001110100111;
		16'b0101001001111110: color_data = 12'b001110100111;
		16'b0101001001111111: color_data = 12'b001110100111;
		16'b0101001010000000: color_data = 12'b001110100111;
		16'b0101001010001101: color_data = 12'b001110100111;
		16'b0101001010001110: color_data = 12'b001110100111;
		16'b0101001010001111: color_data = 12'b001110100111;
		16'b0101001010010000: color_data = 12'b001110100111;
		16'b0101001010010001: color_data = 12'b001110100111;
		16'b0101001010010010: color_data = 12'b001110100111;
		16'b0101001010010011: color_data = 12'b001110100111;
		16'b0101001010010100: color_data = 12'b001110100111;
		16'b0101001010010101: color_data = 12'b001110100111;
		16'b0101001010010110: color_data = 12'b001110100111;
		16'b0101001010010111: color_data = 12'b001110100111;
		16'b0101001010011000: color_data = 12'b001110100111;
		16'b0101001010011001: color_data = 12'b001110100111;
		16'b0101001010100000: color_data = 12'b001110100111;
		16'b0101001010100001: color_data = 12'b001110100111;
		16'b0101001010100010: color_data = 12'b001110100111;
		16'b0101001010100011: color_data = 12'b001110100111;
		16'b0101001010100100: color_data = 12'b001110100111;
		16'b0101001010100101: color_data = 12'b001110100111;
		16'b0101001010100110: color_data = 12'b001110100111;
		16'b0101001010100111: color_data = 12'b001110100111;
		16'b0101001010101000: color_data = 12'b001110100111;
		16'b0101001010101001: color_data = 12'b001110100111;
		16'b0101001010101010: color_data = 12'b001110100111;
		16'b0101001010101011: color_data = 12'b001110100111;
		16'b0101001011001011: color_data = 12'b001110100111;
		16'b0101001011001100: color_data = 12'b001110100111;
		16'b0101001011001101: color_data = 12'b001110100111;
		16'b0101001011001110: color_data = 12'b001110100111;
		16'b0101001011001111: color_data = 12'b001110100111;
		16'b0101001011010000: color_data = 12'b001110100111;
		16'b0101001011010001: color_data = 12'b001110100111;
		16'b0101001011010010: color_data = 12'b001110100111;
		16'b0101001011010011: color_data = 12'b001110100111;
		16'b0101001011010100: color_data = 12'b001110100111;
		16'b0101001011010101: color_data = 12'b001110100111;
		16'b0101001011010110: color_data = 12'b001110100111;
		16'b0101001011010111: color_data = 12'b001110100111;
		16'b0101001011011000: color_data = 12'b001110100111;
		16'b0101001011011001: color_data = 12'b001110100111;
		16'b0101001011011010: color_data = 12'b001110100111;
		16'b0101001011011011: color_data = 12'b001110100111;
		16'b0101001011011100: color_data = 12'b001110100111;
		16'b0101001011011101: color_data = 12'b001110100111;
		16'b0101001011011110: color_data = 12'b001110100111;
		16'b0101001011011111: color_data = 12'b001110100111;
		16'b0101001011100000: color_data = 12'b001110100111;
		16'b0101001011100001: color_data = 12'b001110100111;
		16'b0101001011100010: color_data = 12'b001110100111;
		16'b0101001011100011: color_data = 12'b001110100111;
		16'b0101001011100100: color_data = 12'b001110100111;
		16'b0101001011100101: color_data = 12'b001110100111;
		16'b0101001011100110: color_data = 12'b001110100111;
		16'b0101001011100111: color_data = 12'b001110100111;
		16'b0101001011101000: color_data = 12'b001110100111;
		16'b0101001011110110: color_data = 12'b001110100111;
		16'b0101001011110111: color_data = 12'b001110100111;
		16'b0101001011111000: color_data = 12'b001110100111;
		16'b0101001011111001: color_data = 12'b001110100111;
		16'b0101001011111010: color_data = 12'b001110100111;
		16'b0101001011111011: color_data = 12'b001110100111;
		16'b0101001011111100: color_data = 12'b001110100111;
		16'b0101001011111101: color_data = 12'b001110100111;
		16'b0101001011111110: color_data = 12'b001110100111;
		16'b0101001011111111: color_data = 12'b001110100111;
		16'b0101001100000000: color_data = 12'b001110100111;
		16'b0101001100000001: color_data = 12'b001110100111;
		16'b0101001100011010: color_data = 12'b001110100111;
		16'b0101001100011011: color_data = 12'b001110100111;
		16'b0101001100011100: color_data = 12'b001110100111;
		16'b0101001100011101: color_data = 12'b001110100111;
		16'b0101001100011110: color_data = 12'b001110100111;
		16'b0101001100011111: color_data = 12'b001110100111;
		16'b0101001100100000: color_data = 12'b001110100111;
		16'b0101001100100001: color_data = 12'b001110100111;
		16'b0101001100100010: color_data = 12'b001110100111;
		16'b0101001100100011: color_data = 12'b001110100111;
		16'b0101001100100100: color_data = 12'b001110100111;
		16'b0101001100100101: color_data = 12'b001110100111;
		16'b0101001100100110: color_data = 12'b001110100111;
		16'b0101001100101101: color_data = 12'b001110100111;
		16'b0101001100101110: color_data = 12'b001110100111;
		16'b0101001100101111: color_data = 12'b001110100111;
		16'b0101001100110000: color_data = 12'b001110100111;
		16'b0101001100110001: color_data = 12'b001110100111;
		16'b0101001100110010: color_data = 12'b001110100111;
		16'b0101001100110011: color_data = 12'b001110100111;
		16'b0101001100110100: color_data = 12'b001110100111;
		16'b0101001100110101: color_data = 12'b001110100111;
		16'b0101001100110110: color_data = 12'b001110100111;
		16'b0101001100110111: color_data = 12'b001110100111;
		16'b0101001100111000: color_data = 12'b001110100111;
		16'b0101001101000101: color_data = 12'b001110100111;
		16'b0101001101000110: color_data = 12'b001110100111;
		16'b0101001101000111: color_data = 12'b001110100111;
		16'b0101001101001000: color_data = 12'b001110100111;
		16'b0101001101001001: color_data = 12'b001110100111;
		16'b0101001101001010: color_data = 12'b001110100111;
		16'b0101001101001011: color_data = 12'b001110100111;
		16'b0101001101001100: color_data = 12'b001110100111;
		16'b0101001101001101: color_data = 12'b001110100111;
		16'b0101001101001110: color_data = 12'b001110100111;
		16'b0101001101001111: color_data = 12'b001110100111;
		16'b0101001101010000: color_data = 12'b001110100111;
		16'b0101001101010001: color_data = 12'b001110100111;
		16'b0101001101011000: color_data = 12'b001110100111;
		16'b0101001101011001: color_data = 12'b001110100111;
		16'b0101001101011010: color_data = 12'b001110100111;
		16'b0101001101011011: color_data = 12'b001110100111;
		16'b0101001101011100: color_data = 12'b001110100111;
		16'b0101001101011101: color_data = 12'b001110100111;
		16'b0101001101011110: color_data = 12'b001110100111;
		16'b0101001101011111: color_data = 12'b001110100111;
		16'b0101001101100000: color_data = 12'b001110100111;
		16'b0101001101100001: color_data = 12'b001110100111;
		16'b0101001101100010: color_data = 12'b001110100111;
		16'b0101001101100011: color_data = 12'b001110100111;
		16'b0101010000000000: color_data = 12'b001110100111;
		16'b0101010000000001: color_data = 12'b001110100111;
		16'b0101010000000010: color_data = 12'b001110100111;
		16'b0101010000000011: color_data = 12'b001110100111;
		16'b0101010000000100: color_data = 12'b001110100111;
		16'b0101010000000101: color_data = 12'b001110100111;
		16'b0101010000000110: color_data = 12'b001110100111;
		16'b0101010000000111: color_data = 12'b001110100111;
		16'b0101010000001000: color_data = 12'b001110100111;
		16'b0101010000001001: color_data = 12'b001110100111;
		16'b0101010000001010: color_data = 12'b001110100111;
		16'b0101010000001011: color_data = 12'b001110100111;
		16'b0101010000001100: color_data = 12'b001110100111;
		16'b0101010000101011: color_data = 12'b001110100111;
		16'b0101010000101100: color_data = 12'b001110100111;
		16'b0101010000101101: color_data = 12'b001110100111;
		16'b0101010000101110: color_data = 12'b001110100111;
		16'b0101010000101111: color_data = 12'b001110100111;
		16'b0101010000110000: color_data = 12'b001110100111;
		16'b0101010000110001: color_data = 12'b001110100111;
		16'b0101010000110010: color_data = 12'b001110100111;
		16'b0101010000110011: color_data = 12'b001110100111;
		16'b0101010000110100: color_data = 12'b001110100111;
		16'b0101010000110101: color_data = 12'b001110100111;
		16'b0101010000110110: color_data = 12'b001110100111;
		16'b0101010000110111: color_data = 12'b001110100111;
		16'b0101010000111000: color_data = 12'b001110100111;
		16'b0101010000111001: color_data = 12'b001110100111;
		16'b0101010000111010: color_data = 12'b001110100111;
		16'b0101010000111011: color_data = 12'b001110100111;
		16'b0101010000111100: color_data = 12'b001110100111;
		16'b0101010000111101: color_data = 12'b001110100111;
		16'b0101010000111110: color_data = 12'b001110100111;
		16'b0101010000111111: color_data = 12'b001110100111;
		16'b0101010001000000: color_data = 12'b001110100111;
		16'b0101010001000001: color_data = 12'b001110100111;
		16'b0101010001000010: color_data = 12'b001110100111;
		16'b0101010001000011: color_data = 12'b001110100111;
		16'b0101010001000100: color_data = 12'b001110100111;
		16'b0101010001000101: color_data = 12'b001110100111;
		16'b0101010001000110: color_data = 12'b001110100111;
		16'b0101010001000111: color_data = 12'b001110100111;
		16'b0101010001001000: color_data = 12'b001110100111;
		16'b0101010001001001: color_data = 12'b001110100111;
		16'b0101010001001010: color_data = 12'b001110100111;
		16'b0101010001001011: color_data = 12'b001110100111;
		16'b0101010001001100: color_data = 12'b001110100111;
		16'b0101010001001101: color_data = 12'b001110100111;
		16'b0101010001001110: color_data = 12'b001110100111;
		16'b0101010001001111: color_data = 12'b001110100111;
		16'b0101010001011100: color_data = 12'b001110100111;
		16'b0101010001011101: color_data = 12'b001110100111;
		16'b0101010001011110: color_data = 12'b001110100111;
		16'b0101010001011111: color_data = 12'b001110100111;
		16'b0101010001100000: color_data = 12'b001110100111;
		16'b0101010001100001: color_data = 12'b001110100111;
		16'b0101010001100010: color_data = 12'b001110100111;
		16'b0101010001100011: color_data = 12'b001110100111;
		16'b0101010001100100: color_data = 12'b001110100111;
		16'b0101010001100101: color_data = 12'b001110100111;
		16'b0101010001100110: color_data = 12'b001110100111;
		16'b0101010001100111: color_data = 12'b001110100111;
		16'b0101010001101000: color_data = 12'b001110100111;
		16'b0101010001110101: color_data = 12'b001110100111;
		16'b0101010001110110: color_data = 12'b001110100111;
		16'b0101010001110111: color_data = 12'b001110100111;
		16'b0101010001111000: color_data = 12'b001110100111;
		16'b0101010001111001: color_data = 12'b001110100111;
		16'b0101010001111010: color_data = 12'b001110100111;
		16'b0101010001111011: color_data = 12'b001110100111;
		16'b0101010001111100: color_data = 12'b001110100111;
		16'b0101010001111101: color_data = 12'b001110100111;
		16'b0101010001111110: color_data = 12'b001110100111;
		16'b0101010001111111: color_data = 12'b001110100111;
		16'b0101010010000000: color_data = 12'b001110100111;
		16'b0101010010001101: color_data = 12'b001110100111;
		16'b0101010010001110: color_data = 12'b001110100111;
		16'b0101010010001111: color_data = 12'b001110100111;
		16'b0101010010010000: color_data = 12'b001110100111;
		16'b0101010010010001: color_data = 12'b001110100111;
		16'b0101010010010010: color_data = 12'b001110100111;
		16'b0101010010010011: color_data = 12'b001110100111;
		16'b0101010010010100: color_data = 12'b001110100111;
		16'b0101010010010101: color_data = 12'b001110100111;
		16'b0101010010010110: color_data = 12'b001110100111;
		16'b0101010010010111: color_data = 12'b001110100111;
		16'b0101010010011000: color_data = 12'b001110100111;
		16'b0101010010011001: color_data = 12'b001110100111;
		16'b0101010010100000: color_data = 12'b001110100111;
		16'b0101010010100001: color_data = 12'b001110100111;
		16'b0101010010100010: color_data = 12'b001110100111;
		16'b0101010010100011: color_data = 12'b001110100111;
		16'b0101010010100100: color_data = 12'b001110100111;
		16'b0101010010100101: color_data = 12'b001110100111;
		16'b0101010010100110: color_data = 12'b001110100111;
		16'b0101010010100111: color_data = 12'b001110100111;
		16'b0101010010101000: color_data = 12'b001110100111;
		16'b0101010010101001: color_data = 12'b001110100111;
		16'b0101010010101010: color_data = 12'b001110100111;
		16'b0101010010101011: color_data = 12'b001110100111;
		16'b0101010011001011: color_data = 12'b001110100111;
		16'b0101010011001100: color_data = 12'b001110100111;
		16'b0101010011001101: color_data = 12'b001110100111;
		16'b0101010011001110: color_data = 12'b001110100111;
		16'b0101010011001111: color_data = 12'b001110100111;
		16'b0101010011010000: color_data = 12'b001110100111;
		16'b0101010011010001: color_data = 12'b001110100111;
		16'b0101010011010010: color_data = 12'b001110100111;
		16'b0101010011010011: color_data = 12'b001110100111;
		16'b0101010011010100: color_data = 12'b001110100111;
		16'b0101010011010101: color_data = 12'b001110100111;
		16'b0101010011010110: color_data = 12'b001110100111;
		16'b0101010011010111: color_data = 12'b001110100111;
		16'b0101010011011000: color_data = 12'b001110100111;
		16'b0101010011011001: color_data = 12'b001110100111;
		16'b0101010011011010: color_data = 12'b001110100111;
		16'b0101010011011011: color_data = 12'b001110100111;
		16'b0101010011011100: color_data = 12'b001110100111;
		16'b0101010011011101: color_data = 12'b001110100111;
		16'b0101010011011110: color_data = 12'b001110100111;
		16'b0101010011011111: color_data = 12'b001110100111;
		16'b0101010011100000: color_data = 12'b001110100111;
		16'b0101010011100001: color_data = 12'b001110100111;
		16'b0101010011100010: color_data = 12'b001110100111;
		16'b0101010011100011: color_data = 12'b001110100111;
		16'b0101010011100100: color_data = 12'b001110100111;
		16'b0101010011100101: color_data = 12'b001110100111;
		16'b0101010011100110: color_data = 12'b001110100111;
		16'b0101010011100111: color_data = 12'b001110100111;
		16'b0101010011101000: color_data = 12'b001110100111;
		16'b0101010011110110: color_data = 12'b001110100111;
		16'b0101010011110111: color_data = 12'b001110100111;
		16'b0101010011111000: color_data = 12'b001110100111;
		16'b0101010011111001: color_data = 12'b001110100111;
		16'b0101010011111010: color_data = 12'b001110100111;
		16'b0101010011111011: color_data = 12'b001110100111;
		16'b0101010011111100: color_data = 12'b001110100111;
		16'b0101010011111101: color_data = 12'b001110100111;
		16'b0101010011111110: color_data = 12'b001110100111;
		16'b0101010011111111: color_data = 12'b001110100111;
		16'b0101010100000000: color_data = 12'b001110100111;
		16'b0101010100000001: color_data = 12'b001110100111;
		16'b0101010100011010: color_data = 12'b001110100111;
		16'b0101010100011011: color_data = 12'b001110100111;
		16'b0101010100011100: color_data = 12'b001110100111;
		16'b0101010100011101: color_data = 12'b001110100111;
		16'b0101010100011110: color_data = 12'b001110100111;
		16'b0101010100011111: color_data = 12'b001110100111;
		16'b0101010100100000: color_data = 12'b001110100111;
		16'b0101010100100001: color_data = 12'b001110100111;
		16'b0101010100100010: color_data = 12'b001110100111;
		16'b0101010100100011: color_data = 12'b001110100111;
		16'b0101010100100100: color_data = 12'b001110100111;
		16'b0101010100100101: color_data = 12'b001110100111;
		16'b0101010100100110: color_data = 12'b001110100111;
		16'b0101010100101101: color_data = 12'b001110100111;
		16'b0101010100101110: color_data = 12'b001110100111;
		16'b0101010100101111: color_data = 12'b001110100111;
		16'b0101010100110000: color_data = 12'b001110100111;
		16'b0101010100110001: color_data = 12'b001110100111;
		16'b0101010100110010: color_data = 12'b001110100111;
		16'b0101010100110011: color_data = 12'b001110100111;
		16'b0101010100110100: color_data = 12'b001110100111;
		16'b0101010100110101: color_data = 12'b001110100111;
		16'b0101010100110110: color_data = 12'b001110100111;
		16'b0101010100110111: color_data = 12'b001110100111;
		16'b0101010100111000: color_data = 12'b001110100111;
		16'b0101010101000101: color_data = 12'b001110100111;
		16'b0101010101000110: color_data = 12'b001110100111;
		16'b0101010101000111: color_data = 12'b001110100111;
		16'b0101010101001000: color_data = 12'b001110100111;
		16'b0101010101001001: color_data = 12'b001110100111;
		16'b0101010101001010: color_data = 12'b001110100111;
		16'b0101010101001011: color_data = 12'b001110100111;
		16'b0101010101001100: color_data = 12'b001110100111;
		16'b0101010101001101: color_data = 12'b001110100111;
		16'b0101010101001110: color_data = 12'b001110100111;
		16'b0101010101001111: color_data = 12'b001110100111;
		16'b0101010101010000: color_data = 12'b001110100111;
		16'b0101010101010001: color_data = 12'b001110100111;
		16'b0101010101011000: color_data = 12'b001110100111;
		16'b0101010101011001: color_data = 12'b001110100111;
		16'b0101010101011010: color_data = 12'b001110100111;
		16'b0101010101011011: color_data = 12'b001110100111;
		16'b0101010101011100: color_data = 12'b001110100111;
		16'b0101010101011101: color_data = 12'b001110100111;
		16'b0101010101011110: color_data = 12'b001110100111;
		16'b0101010101011111: color_data = 12'b001110100111;
		16'b0101010101100000: color_data = 12'b001110100111;
		16'b0101010101100001: color_data = 12'b001110100111;
		16'b0101010101100010: color_data = 12'b001110100111;
		16'b0101010101100011: color_data = 12'b001110100111;
		16'b0101011000000000: color_data = 12'b001110100111;
		16'b0101011000000001: color_data = 12'b001110100111;
		16'b0101011000000010: color_data = 12'b001110100111;
		16'b0101011000000011: color_data = 12'b001110100111;
		16'b0101011000000100: color_data = 12'b001110100111;
		16'b0101011000000101: color_data = 12'b001110100111;
		16'b0101011000000110: color_data = 12'b001110100111;
		16'b0101011000000111: color_data = 12'b001110100111;
		16'b0101011000001000: color_data = 12'b001110100111;
		16'b0101011000001001: color_data = 12'b001110100111;
		16'b0101011000001010: color_data = 12'b001110100111;
		16'b0101011000001011: color_data = 12'b001110100111;
		16'b0101011000001100: color_data = 12'b001110100111;
		16'b0101011000101011: color_data = 12'b001110100111;
		16'b0101011000101100: color_data = 12'b001110100111;
		16'b0101011000101101: color_data = 12'b001110100111;
		16'b0101011000101110: color_data = 12'b001110100111;
		16'b0101011000101111: color_data = 12'b001110100111;
		16'b0101011000110000: color_data = 12'b001110100111;
		16'b0101011000110001: color_data = 12'b001110100111;
		16'b0101011000110010: color_data = 12'b001110100111;
		16'b0101011000110011: color_data = 12'b001110100111;
		16'b0101011000110100: color_data = 12'b001110100111;
		16'b0101011000110101: color_data = 12'b001110100111;
		16'b0101011000110110: color_data = 12'b001110100111;
		16'b0101011000110111: color_data = 12'b001110100111;
		16'b0101011000111000: color_data = 12'b001110100111;
		16'b0101011000111001: color_data = 12'b001110100111;
		16'b0101011000111010: color_data = 12'b001110100111;
		16'b0101011000111011: color_data = 12'b001110100111;
		16'b0101011000111100: color_data = 12'b001110100111;
		16'b0101011000111101: color_data = 12'b001110100111;
		16'b0101011000111110: color_data = 12'b001110100111;
		16'b0101011000111111: color_data = 12'b001110100111;
		16'b0101011001000000: color_data = 12'b001110100111;
		16'b0101011001000001: color_data = 12'b001110100111;
		16'b0101011001000010: color_data = 12'b001110100111;
		16'b0101011001000011: color_data = 12'b001110100111;
		16'b0101011001000100: color_data = 12'b001110100111;
		16'b0101011001000101: color_data = 12'b001110100111;
		16'b0101011001000110: color_data = 12'b001110100111;
		16'b0101011001000111: color_data = 12'b001110100111;
		16'b0101011001001000: color_data = 12'b001110100111;
		16'b0101011001001001: color_data = 12'b001110100111;
		16'b0101011001001010: color_data = 12'b001110100111;
		16'b0101011001001011: color_data = 12'b001110100111;
		16'b0101011001001100: color_data = 12'b001110100111;
		16'b0101011001001101: color_data = 12'b001110100111;
		16'b0101011001001110: color_data = 12'b001110100111;
		16'b0101011001001111: color_data = 12'b001110100111;
		16'b0101011001011100: color_data = 12'b001110100111;
		16'b0101011001011101: color_data = 12'b001110100111;
		16'b0101011001011110: color_data = 12'b001110100111;
		16'b0101011001011111: color_data = 12'b001110100111;
		16'b0101011001100000: color_data = 12'b001110100111;
		16'b0101011001100001: color_data = 12'b001110100111;
		16'b0101011001100010: color_data = 12'b001110100111;
		16'b0101011001100011: color_data = 12'b001110100111;
		16'b0101011001100100: color_data = 12'b001110100111;
		16'b0101011001100101: color_data = 12'b001110100111;
		16'b0101011001100110: color_data = 12'b001110100111;
		16'b0101011001100111: color_data = 12'b001110100111;
		16'b0101011001101000: color_data = 12'b001110100111;
		16'b0101011001110101: color_data = 12'b001110100111;
		16'b0101011001110110: color_data = 12'b001110100111;
		16'b0101011001110111: color_data = 12'b001110100111;
		16'b0101011001111000: color_data = 12'b001110100111;
		16'b0101011001111001: color_data = 12'b001110100111;
		16'b0101011001111010: color_data = 12'b001110100111;
		16'b0101011001111011: color_data = 12'b001110100111;
		16'b0101011001111100: color_data = 12'b001110100111;
		16'b0101011001111101: color_data = 12'b001110100111;
		16'b0101011001111110: color_data = 12'b001110100111;
		16'b0101011001111111: color_data = 12'b001110100111;
		16'b0101011010000000: color_data = 12'b001110100111;
		16'b0101011010001101: color_data = 12'b001110100111;
		16'b0101011010001110: color_data = 12'b001110100111;
		16'b0101011010001111: color_data = 12'b001110100111;
		16'b0101011010010000: color_data = 12'b001110100111;
		16'b0101011010010001: color_data = 12'b001110100111;
		16'b0101011010010010: color_data = 12'b001110100111;
		16'b0101011010010011: color_data = 12'b001110100111;
		16'b0101011010010100: color_data = 12'b001110100111;
		16'b0101011010010101: color_data = 12'b001110100111;
		16'b0101011010010110: color_data = 12'b001110100111;
		16'b0101011010010111: color_data = 12'b001110100111;
		16'b0101011010011000: color_data = 12'b001110100111;
		16'b0101011010011001: color_data = 12'b001110100111;
		16'b0101011010100000: color_data = 12'b001110100111;
		16'b0101011010100001: color_data = 12'b001110100111;
		16'b0101011010100010: color_data = 12'b001110100111;
		16'b0101011010100011: color_data = 12'b001110100111;
		16'b0101011010100100: color_data = 12'b001110100111;
		16'b0101011010100101: color_data = 12'b001110100111;
		16'b0101011010100110: color_data = 12'b001110100111;
		16'b0101011010100111: color_data = 12'b001110100111;
		16'b0101011010101000: color_data = 12'b001110100111;
		16'b0101011010101001: color_data = 12'b001110100111;
		16'b0101011010101010: color_data = 12'b001110100111;
		16'b0101011010101011: color_data = 12'b001110100111;
		16'b0101011011001011: color_data = 12'b001110100111;
		16'b0101011011001100: color_data = 12'b001110100111;
		16'b0101011011001101: color_data = 12'b001110100111;
		16'b0101011011001110: color_data = 12'b001110100111;
		16'b0101011011001111: color_data = 12'b001110100111;
		16'b0101011011010000: color_data = 12'b001110100111;
		16'b0101011011010001: color_data = 12'b001110100111;
		16'b0101011011010010: color_data = 12'b001110100111;
		16'b0101011011010011: color_data = 12'b001110100111;
		16'b0101011011010100: color_data = 12'b001110100111;
		16'b0101011011010101: color_data = 12'b001110100111;
		16'b0101011011010110: color_data = 12'b001110100111;
		16'b0101011011010111: color_data = 12'b001110100111;
		16'b0101011011011000: color_data = 12'b001110100111;
		16'b0101011011011001: color_data = 12'b001110100111;
		16'b0101011011011010: color_data = 12'b001110100111;
		16'b0101011011011011: color_data = 12'b001110100111;
		16'b0101011011011100: color_data = 12'b001110100111;
		16'b0101011011011101: color_data = 12'b001110100111;
		16'b0101011011011110: color_data = 12'b001110100111;
		16'b0101011011011111: color_data = 12'b001110100111;
		16'b0101011011100000: color_data = 12'b001110100111;
		16'b0101011011100001: color_data = 12'b001110100111;
		16'b0101011011100010: color_data = 12'b001110100111;
		16'b0101011011100011: color_data = 12'b001110100111;
		16'b0101011011100100: color_data = 12'b001110100111;
		16'b0101011011100101: color_data = 12'b001110100111;
		16'b0101011011100110: color_data = 12'b001110100111;
		16'b0101011011100111: color_data = 12'b001110100111;
		16'b0101011011101000: color_data = 12'b001110100111;
		16'b0101011011110110: color_data = 12'b001110100111;
		16'b0101011011110111: color_data = 12'b001110100111;
		16'b0101011011111000: color_data = 12'b001110100111;
		16'b0101011011111001: color_data = 12'b001110100111;
		16'b0101011011111010: color_data = 12'b001110100111;
		16'b0101011011111011: color_data = 12'b001110100111;
		16'b0101011011111100: color_data = 12'b001110100111;
		16'b0101011011111101: color_data = 12'b001110100111;
		16'b0101011011111110: color_data = 12'b001110100111;
		16'b0101011011111111: color_data = 12'b001110100111;
		16'b0101011100000000: color_data = 12'b001110100111;
		16'b0101011100000001: color_data = 12'b001110100111;
		16'b0101011100011010: color_data = 12'b001110100111;
		16'b0101011100011011: color_data = 12'b001110100111;
		16'b0101011100011100: color_data = 12'b001110100111;
		16'b0101011100011101: color_data = 12'b001110100111;
		16'b0101011100011110: color_data = 12'b001110100111;
		16'b0101011100011111: color_data = 12'b001110100111;
		16'b0101011100100000: color_data = 12'b001110100111;
		16'b0101011100100001: color_data = 12'b001110100111;
		16'b0101011100100010: color_data = 12'b001110100111;
		16'b0101011100100011: color_data = 12'b001110100111;
		16'b0101011100100100: color_data = 12'b001110100111;
		16'b0101011100100101: color_data = 12'b001110100111;
		16'b0101011100100110: color_data = 12'b001110100111;
		16'b0101011100101101: color_data = 12'b001110100111;
		16'b0101011100101110: color_data = 12'b001110100111;
		16'b0101011100101111: color_data = 12'b001110100111;
		16'b0101011100110000: color_data = 12'b001110100111;
		16'b0101011100110001: color_data = 12'b001110100111;
		16'b0101011100110010: color_data = 12'b001110100111;
		16'b0101011100110011: color_data = 12'b001110100111;
		16'b0101011100110100: color_data = 12'b001110100111;
		16'b0101011100110101: color_data = 12'b001110100111;
		16'b0101011100110110: color_data = 12'b001110100111;
		16'b0101011100110111: color_data = 12'b001110100111;
		16'b0101011100111000: color_data = 12'b001110100111;
		16'b0101011101000101: color_data = 12'b001110100111;
		16'b0101011101000110: color_data = 12'b001110100111;
		16'b0101011101000111: color_data = 12'b001110100111;
		16'b0101011101001000: color_data = 12'b001110100111;
		16'b0101011101001001: color_data = 12'b001110100111;
		16'b0101011101001010: color_data = 12'b001110100111;
		16'b0101011101001011: color_data = 12'b001110100111;
		16'b0101011101001100: color_data = 12'b001110100111;
		16'b0101011101001101: color_data = 12'b001110100111;
		16'b0101011101001110: color_data = 12'b001110100111;
		16'b0101011101001111: color_data = 12'b001110100111;
		16'b0101011101010000: color_data = 12'b001110100111;
		16'b0101011101010001: color_data = 12'b001110100111;
		16'b0101011101011000: color_data = 12'b001110100111;
		16'b0101011101011001: color_data = 12'b001110100111;
		16'b0101011101011010: color_data = 12'b001110100111;
		16'b0101011101011011: color_data = 12'b001110100111;
		16'b0101011101011100: color_data = 12'b001110100111;
		16'b0101011101011101: color_data = 12'b001110100111;
		16'b0101011101011110: color_data = 12'b001110100111;
		16'b0101011101011111: color_data = 12'b001110100111;
		16'b0101011101100000: color_data = 12'b001110100111;
		16'b0101011101100001: color_data = 12'b001110100111;
		16'b0101011101100010: color_data = 12'b001110100111;
		16'b0101011101100011: color_data = 12'b001110100111;
		16'b0101100000000000: color_data = 12'b001110100111;
		16'b0101100000000001: color_data = 12'b001110100111;
		16'b0101100000000010: color_data = 12'b001110100111;
		16'b0101100000000011: color_data = 12'b001110100111;
		16'b0101100000000100: color_data = 12'b001110100111;
		16'b0101100000000101: color_data = 12'b001110100111;
		16'b0101100000000110: color_data = 12'b001110100111;
		16'b0101100000000111: color_data = 12'b001110100111;
		16'b0101100000001000: color_data = 12'b001110100111;
		16'b0101100000001001: color_data = 12'b001110100111;
		16'b0101100000001010: color_data = 12'b001110100111;
		16'b0101100000001011: color_data = 12'b001110100111;
		16'b0101100000001100: color_data = 12'b001110100111;
		16'b0101100000101011: color_data = 12'b001110100111;
		16'b0101100000101100: color_data = 12'b001110100111;
		16'b0101100000101101: color_data = 12'b001110100111;
		16'b0101100000101110: color_data = 12'b001110100111;
		16'b0101100000101111: color_data = 12'b001110100111;
		16'b0101100000110000: color_data = 12'b001110100111;
		16'b0101100000110001: color_data = 12'b001110100111;
		16'b0101100000110010: color_data = 12'b001110100111;
		16'b0101100000110011: color_data = 12'b001110100111;
		16'b0101100000110100: color_data = 12'b001110100111;
		16'b0101100000110101: color_data = 12'b001110100111;
		16'b0101100000110110: color_data = 12'b001110100111;
		16'b0101100000110111: color_data = 12'b001110100111;
		16'b0101100000111000: color_data = 12'b001110100111;
		16'b0101100000111001: color_data = 12'b001110100111;
		16'b0101100000111010: color_data = 12'b001110100111;
		16'b0101100000111011: color_data = 12'b001110100111;
		16'b0101100000111100: color_data = 12'b001110100111;
		16'b0101100000111101: color_data = 12'b001110100111;
		16'b0101100000111110: color_data = 12'b001110100111;
		16'b0101100000111111: color_data = 12'b001110100111;
		16'b0101100001000000: color_data = 12'b001110100111;
		16'b0101100001000001: color_data = 12'b001110100111;
		16'b0101100001000010: color_data = 12'b001110100111;
		16'b0101100001000011: color_data = 12'b001110100111;
		16'b0101100001000100: color_data = 12'b001110100111;
		16'b0101100001000101: color_data = 12'b001110100111;
		16'b0101100001000110: color_data = 12'b001110100111;
		16'b0101100001000111: color_data = 12'b001110100111;
		16'b0101100001001000: color_data = 12'b001110100111;
		16'b0101100001001001: color_data = 12'b001110100111;
		16'b0101100001001010: color_data = 12'b001110100111;
		16'b0101100001001011: color_data = 12'b001110100111;
		16'b0101100001001100: color_data = 12'b001110100111;
		16'b0101100001001101: color_data = 12'b001110100111;
		16'b0101100001001110: color_data = 12'b001110100111;
		16'b0101100001001111: color_data = 12'b001110100111;
		16'b0101100001011100: color_data = 12'b001110100111;
		16'b0101100001011101: color_data = 12'b001110100111;
		16'b0101100001011110: color_data = 12'b001110100111;
		16'b0101100001011111: color_data = 12'b001110100111;
		16'b0101100001100000: color_data = 12'b001110100111;
		16'b0101100001100001: color_data = 12'b001110100111;
		16'b0101100001100010: color_data = 12'b001110100111;
		16'b0101100001100011: color_data = 12'b001110100111;
		16'b0101100001100100: color_data = 12'b001110100111;
		16'b0101100001100101: color_data = 12'b001110100111;
		16'b0101100001100110: color_data = 12'b001110100111;
		16'b0101100001100111: color_data = 12'b001110100111;
		16'b0101100001101000: color_data = 12'b001110100111;
		16'b0101100001110101: color_data = 12'b001110100111;
		16'b0101100001110110: color_data = 12'b001110100111;
		16'b0101100001110111: color_data = 12'b001110100111;
		16'b0101100001111000: color_data = 12'b001110100111;
		16'b0101100001111001: color_data = 12'b001110100111;
		16'b0101100001111010: color_data = 12'b001110100111;
		16'b0101100001111011: color_data = 12'b001110100111;
		16'b0101100001111100: color_data = 12'b001110100111;
		16'b0101100001111101: color_data = 12'b001110100111;
		16'b0101100001111110: color_data = 12'b001110100111;
		16'b0101100001111111: color_data = 12'b001110100111;
		16'b0101100010000000: color_data = 12'b001110100111;
		16'b0101100010001101: color_data = 12'b001110100111;
		16'b0101100010001110: color_data = 12'b001110100111;
		16'b0101100010001111: color_data = 12'b001110100111;
		16'b0101100010010000: color_data = 12'b001110100111;
		16'b0101100010010001: color_data = 12'b001110100111;
		16'b0101100010010010: color_data = 12'b001110100111;
		16'b0101100010010011: color_data = 12'b001110100111;
		16'b0101100010010100: color_data = 12'b001110100111;
		16'b0101100010010101: color_data = 12'b001110100111;
		16'b0101100010010110: color_data = 12'b001110100111;
		16'b0101100010010111: color_data = 12'b001110100111;
		16'b0101100010011000: color_data = 12'b001110100111;
		16'b0101100010011001: color_data = 12'b001110100111;
		16'b0101100010100000: color_data = 12'b001110100111;
		16'b0101100010100001: color_data = 12'b001110100111;
		16'b0101100010100010: color_data = 12'b001110100111;
		16'b0101100010100011: color_data = 12'b001110100111;
		16'b0101100010100100: color_data = 12'b001110100111;
		16'b0101100010100101: color_data = 12'b001110100111;
		16'b0101100010100110: color_data = 12'b001110100111;
		16'b0101100010100111: color_data = 12'b001110100111;
		16'b0101100010101000: color_data = 12'b001110100111;
		16'b0101100010101001: color_data = 12'b001110100111;
		16'b0101100010101010: color_data = 12'b001110100111;
		16'b0101100010101011: color_data = 12'b001110100111;
		16'b0101100011001011: color_data = 12'b001110100111;
		16'b0101100011001100: color_data = 12'b001110100111;
		16'b0101100011001101: color_data = 12'b001110100111;
		16'b0101100011001110: color_data = 12'b001110100111;
		16'b0101100011001111: color_data = 12'b001110100111;
		16'b0101100011010000: color_data = 12'b001110100111;
		16'b0101100011010001: color_data = 12'b001110100111;
		16'b0101100011010010: color_data = 12'b001110100111;
		16'b0101100011010011: color_data = 12'b001110100111;
		16'b0101100011010100: color_data = 12'b001110100111;
		16'b0101100011010101: color_data = 12'b001110100111;
		16'b0101100011010110: color_data = 12'b001110100111;
		16'b0101100011010111: color_data = 12'b001110100111;
		16'b0101100011011000: color_data = 12'b001110100111;
		16'b0101100011011001: color_data = 12'b001110100111;
		16'b0101100011011010: color_data = 12'b001110100111;
		16'b0101100011011011: color_data = 12'b001110100111;
		16'b0101100011011100: color_data = 12'b001110100111;
		16'b0101100011011101: color_data = 12'b001110100111;
		16'b0101100011011110: color_data = 12'b001110100111;
		16'b0101100011011111: color_data = 12'b001110100111;
		16'b0101100011100000: color_data = 12'b001110100111;
		16'b0101100011100001: color_data = 12'b001110100111;
		16'b0101100011100010: color_data = 12'b001110100111;
		16'b0101100011100011: color_data = 12'b001110100111;
		16'b0101100011100100: color_data = 12'b001110100111;
		16'b0101100011100101: color_data = 12'b001110100111;
		16'b0101100011100110: color_data = 12'b001110100111;
		16'b0101100011100111: color_data = 12'b001110100111;
		16'b0101100011101000: color_data = 12'b001110100111;
		16'b0101100011110110: color_data = 12'b001110100111;
		16'b0101100011110111: color_data = 12'b001110100111;
		16'b0101100011111000: color_data = 12'b001110100111;
		16'b0101100011111001: color_data = 12'b001110100111;
		16'b0101100011111010: color_data = 12'b001110100111;
		16'b0101100011111011: color_data = 12'b001110100111;
		16'b0101100011111100: color_data = 12'b001110100111;
		16'b0101100011111101: color_data = 12'b001110100111;
		16'b0101100011111110: color_data = 12'b001110100111;
		16'b0101100011111111: color_data = 12'b001110100111;
		16'b0101100100000000: color_data = 12'b001110100111;
		16'b0101100100000001: color_data = 12'b001110100111;
		16'b0101100100011010: color_data = 12'b001110100111;
		16'b0101100100011011: color_data = 12'b001110100111;
		16'b0101100100011100: color_data = 12'b001110100111;
		16'b0101100100011101: color_data = 12'b001110100111;
		16'b0101100100011110: color_data = 12'b001110100111;
		16'b0101100100011111: color_data = 12'b001110100111;
		16'b0101100100100000: color_data = 12'b001110100111;
		16'b0101100100100001: color_data = 12'b001110100111;
		16'b0101100100100010: color_data = 12'b001110100111;
		16'b0101100100100011: color_data = 12'b001110100111;
		16'b0101100100100100: color_data = 12'b001110100111;
		16'b0101100100100101: color_data = 12'b001110100111;
		16'b0101100100100110: color_data = 12'b001110100111;
		16'b0101100100101101: color_data = 12'b001110100111;
		16'b0101100100101110: color_data = 12'b001110100111;
		16'b0101100100101111: color_data = 12'b001110100111;
		16'b0101100100110000: color_data = 12'b001110100111;
		16'b0101100100110001: color_data = 12'b001110100111;
		16'b0101100100110010: color_data = 12'b001110100111;
		16'b0101100100110011: color_data = 12'b001110100111;
		16'b0101100100110100: color_data = 12'b001110100111;
		16'b0101100100110101: color_data = 12'b001110100111;
		16'b0101100100110110: color_data = 12'b001110100111;
		16'b0101100100110111: color_data = 12'b001110100111;
		16'b0101100100111000: color_data = 12'b001110100111;
		16'b0101100101000101: color_data = 12'b001110100111;
		16'b0101100101000110: color_data = 12'b001110100111;
		16'b0101100101000111: color_data = 12'b001110100111;
		16'b0101100101001000: color_data = 12'b001110100111;
		16'b0101100101001001: color_data = 12'b001110100111;
		16'b0101100101001010: color_data = 12'b001110100111;
		16'b0101100101001011: color_data = 12'b001110100111;
		16'b0101100101001100: color_data = 12'b001110100111;
		16'b0101100101001101: color_data = 12'b001110100111;
		16'b0101100101001110: color_data = 12'b001110100111;
		16'b0101100101001111: color_data = 12'b001110100111;
		16'b0101100101010000: color_data = 12'b001110100111;
		16'b0101100101010001: color_data = 12'b001110100111;
		16'b0101100101011000: color_data = 12'b001110100111;
		16'b0101100101011001: color_data = 12'b001110100111;
		16'b0101100101011010: color_data = 12'b001110100111;
		16'b0101100101011011: color_data = 12'b001110100111;
		16'b0101100101011100: color_data = 12'b001110100111;
		16'b0101100101011101: color_data = 12'b001110100111;
		16'b0101100101011110: color_data = 12'b001110100111;
		16'b0101100101011111: color_data = 12'b001110100111;
		16'b0101100101100000: color_data = 12'b001110100111;
		16'b0101100101100001: color_data = 12'b001110100111;
		16'b0101100101100010: color_data = 12'b001110100111;
		16'b0101100101100011: color_data = 12'b001110100111;
		16'b0101101000000000: color_data = 12'b001110100111;
		16'b0101101000000001: color_data = 12'b001110100111;
		16'b0101101000000010: color_data = 12'b001110100111;
		16'b0101101000000011: color_data = 12'b001110100111;
		16'b0101101000000100: color_data = 12'b001110100111;
		16'b0101101000000101: color_data = 12'b001110100111;
		16'b0101101000000110: color_data = 12'b001110100111;
		16'b0101101000000111: color_data = 12'b001110100111;
		16'b0101101000001000: color_data = 12'b001110100111;
		16'b0101101000001001: color_data = 12'b001110100111;
		16'b0101101000001010: color_data = 12'b001110100111;
		16'b0101101000001011: color_data = 12'b001110100111;
		16'b0101101000001100: color_data = 12'b001110100111;
		16'b0101101000101011: color_data = 12'b001110100111;
		16'b0101101000101100: color_data = 12'b001110100111;
		16'b0101101000101101: color_data = 12'b001110100111;
		16'b0101101000101110: color_data = 12'b001110100111;
		16'b0101101000101111: color_data = 12'b001110100111;
		16'b0101101000110000: color_data = 12'b001110100111;
		16'b0101101000110001: color_data = 12'b001110100111;
		16'b0101101000110010: color_data = 12'b001110100111;
		16'b0101101000110011: color_data = 12'b001110100111;
		16'b0101101000110100: color_data = 12'b001110100111;
		16'b0101101000110101: color_data = 12'b001110100111;
		16'b0101101000110110: color_data = 12'b001110100111;
		16'b0101101000110111: color_data = 12'b001110100111;
		16'b0101101000111000: color_data = 12'b001110100111;
		16'b0101101000111001: color_data = 12'b001110100111;
		16'b0101101000111010: color_data = 12'b001110100111;
		16'b0101101000111011: color_data = 12'b001110100111;
		16'b0101101000111100: color_data = 12'b001110100111;
		16'b0101101000111101: color_data = 12'b001110100111;
		16'b0101101000111110: color_data = 12'b001110100111;
		16'b0101101000111111: color_data = 12'b001110100111;
		16'b0101101001000000: color_data = 12'b001110100111;
		16'b0101101001000001: color_data = 12'b001110100111;
		16'b0101101001000010: color_data = 12'b001110100111;
		16'b0101101001000011: color_data = 12'b001110100111;
		16'b0101101001000100: color_data = 12'b001110100111;
		16'b0101101001000101: color_data = 12'b001110100111;
		16'b0101101001000110: color_data = 12'b001110100111;
		16'b0101101001000111: color_data = 12'b001110100111;
		16'b0101101001001000: color_data = 12'b001110100111;
		16'b0101101001001001: color_data = 12'b001110100111;
		16'b0101101001001010: color_data = 12'b001110100111;
		16'b0101101001001011: color_data = 12'b001110100111;
		16'b0101101001001100: color_data = 12'b001110100111;
		16'b0101101001001101: color_data = 12'b001110100111;
		16'b0101101001001110: color_data = 12'b001110100111;
		16'b0101101001001111: color_data = 12'b001110100111;
		16'b0101101001011100: color_data = 12'b001110100111;
		16'b0101101001011101: color_data = 12'b001110100111;
		16'b0101101001011110: color_data = 12'b001110100111;
		16'b0101101001011111: color_data = 12'b001110100111;
		16'b0101101001100000: color_data = 12'b001110100111;
		16'b0101101001100001: color_data = 12'b001110100111;
		16'b0101101001100010: color_data = 12'b001110100111;
		16'b0101101001100011: color_data = 12'b001110100111;
		16'b0101101001100100: color_data = 12'b001110100111;
		16'b0101101001100101: color_data = 12'b001110100111;
		16'b0101101001100110: color_data = 12'b001110100111;
		16'b0101101001100111: color_data = 12'b001110100111;
		16'b0101101001101000: color_data = 12'b001110100111;
		16'b0101101001110101: color_data = 12'b001110100111;
		16'b0101101001110110: color_data = 12'b001110100111;
		16'b0101101001110111: color_data = 12'b001110100111;
		16'b0101101001111000: color_data = 12'b001110100111;
		16'b0101101001111001: color_data = 12'b001110100111;
		16'b0101101001111010: color_data = 12'b001110100111;
		16'b0101101001111011: color_data = 12'b001110100111;
		16'b0101101001111100: color_data = 12'b001110100111;
		16'b0101101001111101: color_data = 12'b001110100111;
		16'b0101101001111110: color_data = 12'b001110100111;
		16'b0101101001111111: color_data = 12'b001110100111;
		16'b0101101010000000: color_data = 12'b001110100111;
		16'b0101101010001101: color_data = 12'b001110100111;
		16'b0101101010001110: color_data = 12'b001110100111;
		16'b0101101010001111: color_data = 12'b001110100111;
		16'b0101101010010000: color_data = 12'b001110100111;
		16'b0101101010010001: color_data = 12'b001110100111;
		16'b0101101010010010: color_data = 12'b001110100111;
		16'b0101101010010011: color_data = 12'b001110100111;
		16'b0101101010010100: color_data = 12'b001110100111;
		16'b0101101010010101: color_data = 12'b001110100111;
		16'b0101101010010110: color_data = 12'b001110100111;
		16'b0101101010010111: color_data = 12'b001110100111;
		16'b0101101010011000: color_data = 12'b001110100111;
		16'b0101101010011001: color_data = 12'b001110100111;
		16'b0101101010100000: color_data = 12'b001110100111;
		16'b0101101010100001: color_data = 12'b001110100111;
		16'b0101101010100010: color_data = 12'b001110100111;
		16'b0101101010100011: color_data = 12'b001110100111;
		16'b0101101010100100: color_data = 12'b001110100111;
		16'b0101101010100101: color_data = 12'b001110100111;
		16'b0101101010100110: color_data = 12'b001110100111;
		16'b0101101010100111: color_data = 12'b001110100111;
		16'b0101101010101000: color_data = 12'b001110100111;
		16'b0101101010101001: color_data = 12'b001110100111;
		16'b0101101010101010: color_data = 12'b001110100111;
		16'b0101101010101011: color_data = 12'b001110100111;
		16'b0101101011001011: color_data = 12'b001110100111;
		16'b0101101011001100: color_data = 12'b001110100111;
		16'b0101101011001101: color_data = 12'b001110100111;
		16'b0101101011001110: color_data = 12'b001110100111;
		16'b0101101011001111: color_data = 12'b001110100111;
		16'b0101101011010000: color_data = 12'b001110100111;
		16'b0101101011010001: color_data = 12'b001110100111;
		16'b0101101011010010: color_data = 12'b001110100111;
		16'b0101101011010011: color_data = 12'b001110100111;
		16'b0101101011010100: color_data = 12'b001110100111;
		16'b0101101011010101: color_data = 12'b001110100111;
		16'b0101101011010110: color_data = 12'b001110100111;
		16'b0101101011010111: color_data = 12'b001110100111;
		16'b0101101011011000: color_data = 12'b001110100111;
		16'b0101101011011001: color_data = 12'b001110100111;
		16'b0101101011011010: color_data = 12'b001110100111;
		16'b0101101011011011: color_data = 12'b001110100111;
		16'b0101101011011100: color_data = 12'b001110100111;
		16'b0101101011011101: color_data = 12'b001110100111;
		16'b0101101011011110: color_data = 12'b001110100111;
		16'b0101101011011111: color_data = 12'b001110100111;
		16'b0101101011100000: color_data = 12'b001110100111;
		16'b0101101011100001: color_data = 12'b001110100111;
		16'b0101101011100010: color_data = 12'b001110100111;
		16'b0101101011100011: color_data = 12'b001110100111;
		16'b0101101011100100: color_data = 12'b001110100111;
		16'b0101101011100101: color_data = 12'b001110100111;
		16'b0101101011100110: color_data = 12'b001110100111;
		16'b0101101011100111: color_data = 12'b001110100111;
		16'b0101101011101000: color_data = 12'b001110100111;
		16'b0101101011110110: color_data = 12'b001110100111;
		16'b0101101011110111: color_data = 12'b001110100111;
		16'b0101101011111000: color_data = 12'b001110100111;
		16'b0101101011111001: color_data = 12'b001110100111;
		16'b0101101011111010: color_data = 12'b001110100111;
		16'b0101101011111011: color_data = 12'b001110100111;
		16'b0101101011111100: color_data = 12'b001110100111;
		16'b0101101011111101: color_data = 12'b001110100111;
		16'b0101101011111110: color_data = 12'b001110100111;
		16'b0101101011111111: color_data = 12'b001110100111;
		16'b0101101100000000: color_data = 12'b001110100111;
		16'b0101101100000001: color_data = 12'b001110100111;
		16'b0101101100011010: color_data = 12'b001110100111;
		16'b0101101100011011: color_data = 12'b001110100111;
		16'b0101101100011100: color_data = 12'b001110100111;
		16'b0101101100011101: color_data = 12'b001110100111;
		16'b0101101100011110: color_data = 12'b001110100111;
		16'b0101101100011111: color_data = 12'b001110100111;
		16'b0101101100100000: color_data = 12'b001110100111;
		16'b0101101100100001: color_data = 12'b001110100111;
		16'b0101101100100010: color_data = 12'b001110100111;
		16'b0101101100100011: color_data = 12'b001110100111;
		16'b0101101100100100: color_data = 12'b001110100111;
		16'b0101101100100101: color_data = 12'b001110100111;
		16'b0101101100100110: color_data = 12'b001110100111;
		16'b0101101100101101: color_data = 12'b001110100111;
		16'b0101101100101110: color_data = 12'b001110100111;
		16'b0101101100101111: color_data = 12'b001110100111;
		16'b0101101100110000: color_data = 12'b001110100111;
		16'b0101101100110001: color_data = 12'b001110100111;
		16'b0101101100110010: color_data = 12'b001110100111;
		16'b0101101100110011: color_data = 12'b001110100111;
		16'b0101101100110100: color_data = 12'b001110100111;
		16'b0101101100110101: color_data = 12'b001110100111;
		16'b0101101100110110: color_data = 12'b001110100111;
		16'b0101101100110111: color_data = 12'b001110100111;
		16'b0101101100111000: color_data = 12'b001110100111;
		16'b0101101101000101: color_data = 12'b001110100111;
		16'b0101101101000110: color_data = 12'b001110100111;
		16'b0101101101000111: color_data = 12'b001110100111;
		16'b0101101101001000: color_data = 12'b001110100111;
		16'b0101101101001001: color_data = 12'b001110100111;
		16'b0101101101001010: color_data = 12'b001110100111;
		16'b0101101101001011: color_data = 12'b001110100111;
		16'b0101101101001100: color_data = 12'b001110100111;
		16'b0101101101001101: color_data = 12'b001110100111;
		16'b0101101101001110: color_data = 12'b001110100111;
		16'b0101101101001111: color_data = 12'b001110100111;
		16'b0101101101010000: color_data = 12'b001110100111;
		16'b0101101101010001: color_data = 12'b001110100111;
		16'b0101101101011000: color_data = 12'b001110100111;
		16'b0101101101011001: color_data = 12'b001110100111;
		16'b0101101101011010: color_data = 12'b001110100111;
		16'b0101101101011011: color_data = 12'b001110100111;
		16'b0101101101011100: color_data = 12'b001110100111;
		16'b0101101101011101: color_data = 12'b001110100111;
		16'b0101101101011110: color_data = 12'b001110100111;
		16'b0101101101011111: color_data = 12'b001110100111;
		16'b0101101101100000: color_data = 12'b001110100111;
		16'b0101101101100001: color_data = 12'b001110100111;
		16'b0101101101100010: color_data = 12'b001110100111;
		16'b0101101101100011: color_data = 12'b001110100111;
		16'b0101110000000000: color_data = 12'b001110100111;
		16'b0101110000000001: color_data = 12'b001110100111;
		16'b0101110000000010: color_data = 12'b001110100111;
		16'b0101110000000011: color_data = 12'b001110100111;
		16'b0101110000000100: color_data = 12'b001110100111;
		16'b0101110000000101: color_data = 12'b001110100111;
		16'b0101110000000110: color_data = 12'b001110100111;
		16'b0101110000000111: color_data = 12'b001110100111;
		16'b0101110000001000: color_data = 12'b001110100111;
		16'b0101110000001001: color_data = 12'b001110100111;
		16'b0101110000001010: color_data = 12'b001110100111;
		16'b0101110000001011: color_data = 12'b001110100111;
		16'b0101110000001100: color_data = 12'b001110100111;
		16'b0101110000101011: color_data = 12'b001110100111;
		16'b0101110000101100: color_data = 12'b001110100111;
		16'b0101110000101101: color_data = 12'b001110100111;
		16'b0101110000101110: color_data = 12'b001110100111;
		16'b0101110000101111: color_data = 12'b001110100111;
		16'b0101110000110000: color_data = 12'b001110100111;
		16'b0101110000110001: color_data = 12'b001110100111;
		16'b0101110000110010: color_data = 12'b001110100111;
		16'b0101110000110011: color_data = 12'b001110100111;
		16'b0101110000110100: color_data = 12'b001110100111;
		16'b0101110000110101: color_data = 12'b001110100111;
		16'b0101110000110110: color_data = 12'b001110100111;
		16'b0101110000110111: color_data = 12'b001110100111;
		16'b0101110000111000: color_data = 12'b001110100111;
		16'b0101110000111001: color_data = 12'b001110100111;
		16'b0101110000111010: color_data = 12'b001110100111;
		16'b0101110000111011: color_data = 12'b001110100111;
		16'b0101110000111100: color_data = 12'b001110100111;
		16'b0101110000111101: color_data = 12'b001110100111;
		16'b0101110000111110: color_data = 12'b001110100111;
		16'b0101110000111111: color_data = 12'b001110100111;
		16'b0101110001000000: color_data = 12'b001110100111;
		16'b0101110001000001: color_data = 12'b001110100111;
		16'b0101110001000010: color_data = 12'b001110100111;
		16'b0101110001000011: color_data = 12'b001110100111;
		16'b0101110001000100: color_data = 12'b001110100111;
		16'b0101110001000101: color_data = 12'b001110100111;
		16'b0101110001000110: color_data = 12'b001110100111;
		16'b0101110001000111: color_data = 12'b001110100111;
		16'b0101110001001000: color_data = 12'b001110100111;
		16'b0101110001001001: color_data = 12'b001110100111;
		16'b0101110001001010: color_data = 12'b001110100111;
		16'b0101110001001011: color_data = 12'b001110100111;
		16'b0101110001001100: color_data = 12'b001110100111;
		16'b0101110001001101: color_data = 12'b001110100111;
		16'b0101110001001110: color_data = 12'b001110100111;
		16'b0101110001001111: color_data = 12'b001110100111;
		16'b0101110001011100: color_data = 12'b001110100111;
		16'b0101110001011101: color_data = 12'b001110100111;
		16'b0101110001011110: color_data = 12'b001110100111;
		16'b0101110001011111: color_data = 12'b001110100111;
		16'b0101110001100000: color_data = 12'b001110100111;
		16'b0101110001100001: color_data = 12'b001110100111;
		16'b0101110001100010: color_data = 12'b001110100111;
		16'b0101110001100011: color_data = 12'b001110100111;
		16'b0101110001100100: color_data = 12'b001110100111;
		16'b0101110001100101: color_data = 12'b001110100111;
		16'b0101110001100110: color_data = 12'b001110100111;
		16'b0101110001100111: color_data = 12'b001110100111;
		16'b0101110001101000: color_data = 12'b001110100111;
		16'b0101110001110101: color_data = 12'b001110100111;
		16'b0101110001110110: color_data = 12'b001110100111;
		16'b0101110001110111: color_data = 12'b001110100111;
		16'b0101110001111000: color_data = 12'b001110100111;
		16'b0101110001111001: color_data = 12'b001110100111;
		16'b0101110001111010: color_data = 12'b001110100111;
		16'b0101110001111011: color_data = 12'b001110100111;
		16'b0101110001111100: color_data = 12'b001110100111;
		16'b0101110001111101: color_data = 12'b001110100111;
		16'b0101110001111110: color_data = 12'b001110100111;
		16'b0101110001111111: color_data = 12'b001110100111;
		16'b0101110010000000: color_data = 12'b001110100111;
		16'b0101110010001101: color_data = 12'b001110100111;
		16'b0101110010001110: color_data = 12'b001110100111;
		16'b0101110010001111: color_data = 12'b001110100111;
		16'b0101110010010000: color_data = 12'b001110100111;
		16'b0101110010010001: color_data = 12'b001110100111;
		16'b0101110010010010: color_data = 12'b001110100111;
		16'b0101110010010011: color_data = 12'b001110100111;
		16'b0101110010010100: color_data = 12'b001110100111;
		16'b0101110010010101: color_data = 12'b001110100111;
		16'b0101110010010110: color_data = 12'b001110100111;
		16'b0101110010010111: color_data = 12'b001110100111;
		16'b0101110010011000: color_data = 12'b001110100111;
		16'b0101110010011001: color_data = 12'b001110100111;
		16'b0101110010100000: color_data = 12'b001110100111;
		16'b0101110010100001: color_data = 12'b001110100111;
		16'b0101110010100010: color_data = 12'b001110100111;
		16'b0101110010100011: color_data = 12'b001110100111;
		16'b0101110010100100: color_data = 12'b001110100111;
		16'b0101110010100101: color_data = 12'b001110100111;
		16'b0101110010100110: color_data = 12'b001110100111;
		16'b0101110010100111: color_data = 12'b001110100111;
		16'b0101110010101000: color_data = 12'b001110100111;
		16'b0101110010101001: color_data = 12'b001110100111;
		16'b0101110010101010: color_data = 12'b001110100111;
		16'b0101110010101011: color_data = 12'b001110100111;
		16'b0101110011001011: color_data = 12'b001110100111;
		16'b0101110011001100: color_data = 12'b001110100111;
		16'b0101110011001101: color_data = 12'b001110100111;
		16'b0101110011001110: color_data = 12'b001110100111;
		16'b0101110011001111: color_data = 12'b001110100111;
		16'b0101110011010000: color_data = 12'b001110100111;
		16'b0101110011010001: color_data = 12'b001110100111;
		16'b0101110011010010: color_data = 12'b001110100111;
		16'b0101110011010011: color_data = 12'b001110100111;
		16'b0101110011010100: color_data = 12'b001110100111;
		16'b0101110011010101: color_data = 12'b001110100111;
		16'b0101110011010110: color_data = 12'b001110100111;
		16'b0101110011010111: color_data = 12'b001110100111;
		16'b0101110011011000: color_data = 12'b001110100111;
		16'b0101110011011001: color_data = 12'b001110100111;
		16'b0101110011011010: color_data = 12'b001110100111;
		16'b0101110011011011: color_data = 12'b001110100111;
		16'b0101110011011100: color_data = 12'b001110100111;
		16'b0101110011011101: color_data = 12'b001110100111;
		16'b0101110011011110: color_data = 12'b001110100111;
		16'b0101110011011111: color_data = 12'b001110100111;
		16'b0101110011100000: color_data = 12'b001110100111;
		16'b0101110011100001: color_data = 12'b001110100111;
		16'b0101110011100010: color_data = 12'b001110100111;
		16'b0101110011100011: color_data = 12'b001110100111;
		16'b0101110011100100: color_data = 12'b001110100111;
		16'b0101110011100101: color_data = 12'b001110100111;
		16'b0101110011100110: color_data = 12'b001110100111;
		16'b0101110011100111: color_data = 12'b001110100111;
		16'b0101110011101000: color_data = 12'b001110100111;
		16'b0101110011110110: color_data = 12'b001110100111;
		16'b0101110011110111: color_data = 12'b001110100111;
		16'b0101110011111000: color_data = 12'b001110100111;
		16'b0101110011111001: color_data = 12'b001110100111;
		16'b0101110011111010: color_data = 12'b001110100111;
		16'b0101110011111011: color_data = 12'b001110100111;
		16'b0101110011111100: color_data = 12'b001110100111;
		16'b0101110011111101: color_data = 12'b001110100111;
		16'b0101110011111110: color_data = 12'b001110100111;
		16'b0101110011111111: color_data = 12'b001110100111;
		16'b0101110100000000: color_data = 12'b001110100111;
		16'b0101110100000001: color_data = 12'b001110100111;
		16'b0101110100011010: color_data = 12'b001110100111;
		16'b0101110100011011: color_data = 12'b001110100111;
		16'b0101110100011100: color_data = 12'b001110100111;
		16'b0101110100011101: color_data = 12'b001110100111;
		16'b0101110100011110: color_data = 12'b001110100111;
		16'b0101110100011111: color_data = 12'b001110100111;
		16'b0101110100100000: color_data = 12'b001110100111;
		16'b0101110100100001: color_data = 12'b001110100111;
		16'b0101110100100010: color_data = 12'b001110100111;
		16'b0101110100100011: color_data = 12'b001110100111;
		16'b0101110100100100: color_data = 12'b001110100111;
		16'b0101110100100101: color_data = 12'b001110100111;
		16'b0101110100100110: color_data = 12'b001110100111;
		16'b0101110100101101: color_data = 12'b001110100111;
		16'b0101110100101110: color_data = 12'b001110100111;
		16'b0101110100101111: color_data = 12'b001110100111;
		16'b0101110100110000: color_data = 12'b001110100111;
		16'b0101110100110001: color_data = 12'b001110100111;
		16'b0101110100110010: color_data = 12'b001110100111;
		16'b0101110100110011: color_data = 12'b001110100111;
		16'b0101110100110100: color_data = 12'b001110100111;
		16'b0101110100110101: color_data = 12'b001110100111;
		16'b0101110100110110: color_data = 12'b001110100111;
		16'b0101110100110111: color_data = 12'b001110100111;
		16'b0101110100111000: color_data = 12'b001110100111;
		16'b0101110101000101: color_data = 12'b001110100111;
		16'b0101110101000110: color_data = 12'b001110100111;
		16'b0101110101000111: color_data = 12'b001110100111;
		16'b0101110101001000: color_data = 12'b001110100111;
		16'b0101110101001001: color_data = 12'b001110100111;
		16'b0101110101001010: color_data = 12'b001110100111;
		16'b0101110101001011: color_data = 12'b001110100111;
		16'b0101110101001100: color_data = 12'b001110100111;
		16'b0101110101001101: color_data = 12'b001110100111;
		16'b0101110101001110: color_data = 12'b001110100111;
		16'b0101110101001111: color_data = 12'b001110100111;
		16'b0101110101010000: color_data = 12'b001110100111;
		16'b0101110101010001: color_data = 12'b001110100111;
		16'b0101110101011000: color_data = 12'b001110100111;
		16'b0101110101011001: color_data = 12'b001110100111;
		16'b0101110101011010: color_data = 12'b001110100111;
		16'b0101110101011011: color_data = 12'b001110100111;
		16'b0101110101011100: color_data = 12'b001110100111;
		16'b0101110101011101: color_data = 12'b001110100111;
		16'b0101110101011110: color_data = 12'b001110100111;
		16'b0101110101011111: color_data = 12'b001110100111;
		16'b0101110101100000: color_data = 12'b001110100111;
		16'b0101110101100001: color_data = 12'b001110100111;
		16'b0101110101100010: color_data = 12'b001110100111;
		16'b0101110101100011: color_data = 12'b001110100111;
		16'b0101111000000000: color_data = 12'b001110100111;
		16'b0101111000000001: color_data = 12'b001110100111;
		16'b0101111000000010: color_data = 12'b001110100111;
		16'b0101111000000011: color_data = 12'b001110100111;
		16'b0101111000000100: color_data = 12'b001110100111;
		16'b0101111000000101: color_data = 12'b001110100111;
		16'b0101111000000110: color_data = 12'b001110100111;
		16'b0101111000000111: color_data = 12'b001110100111;
		16'b0101111000001000: color_data = 12'b001110100111;
		16'b0101111000001001: color_data = 12'b001110100111;
		16'b0101111000001010: color_data = 12'b001110100111;
		16'b0101111000001011: color_data = 12'b001110100111;
		16'b0101111000001100: color_data = 12'b001110100111;
		16'b0101111000101011: color_data = 12'b001110100111;
		16'b0101111000101100: color_data = 12'b001110100111;
		16'b0101111000101101: color_data = 12'b001110100111;
		16'b0101111000101110: color_data = 12'b001110100111;
		16'b0101111000101111: color_data = 12'b001110100111;
		16'b0101111000110000: color_data = 12'b001110100111;
		16'b0101111000110001: color_data = 12'b001110100111;
		16'b0101111000110010: color_data = 12'b001110100111;
		16'b0101111000110011: color_data = 12'b001110100111;
		16'b0101111000110100: color_data = 12'b001110100111;
		16'b0101111000110101: color_data = 12'b001110100111;
		16'b0101111000110110: color_data = 12'b001110100111;
		16'b0101111000110111: color_data = 12'b001110100111;
		16'b0101111000111000: color_data = 12'b001110100111;
		16'b0101111000111001: color_data = 12'b001110100111;
		16'b0101111000111010: color_data = 12'b001110100111;
		16'b0101111000111011: color_data = 12'b001110100111;
		16'b0101111000111100: color_data = 12'b001110100111;
		16'b0101111000111101: color_data = 12'b001110100111;
		16'b0101111000111110: color_data = 12'b001110100111;
		16'b0101111000111111: color_data = 12'b001110100111;
		16'b0101111001000000: color_data = 12'b001110100111;
		16'b0101111001000001: color_data = 12'b001110100111;
		16'b0101111001000010: color_data = 12'b001110100111;
		16'b0101111001000011: color_data = 12'b001110100111;
		16'b0101111001000100: color_data = 12'b001110100111;
		16'b0101111001000101: color_data = 12'b001110100111;
		16'b0101111001000110: color_data = 12'b001110100111;
		16'b0101111001000111: color_data = 12'b001110100111;
		16'b0101111001001000: color_data = 12'b001110100111;
		16'b0101111001001001: color_data = 12'b001110100111;
		16'b0101111001001010: color_data = 12'b001110100111;
		16'b0101111001001011: color_data = 12'b001110100111;
		16'b0101111001001100: color_data = 12'b001110100111;
		16'b0101111001001101: color_data = 12'b001110100111;
		16'b0101111001001110: color_data = 12'b001110100111;
		16'b0101111001001111: color_data = 12'b001110100111;
		16'b0101111001011100: color_data = 12'b001110100111;
		16'b0101111001011101: color_data = 12'b001110100111;
		16'b0101111001011110: color_data = 12'b001110100111;
		16'b0101111001011111: color_data = 12'b001110100111;
		16'b0101111001100000: color_data = 12'b001110100111;
		16'b0101111001100001: color_data = 12'b001110100111;
		16'b0101111001100010: color_data = 12'b001110100111;
		16'b0101111001100011: color_data = 12'b001110100111;
		16'b0101111001100100: color_data = 12'b001110100111;
		16'b0101111001100101: color_data = 12'b001110100111;
		16'b0101111001100110: color_data = 12'b001110100111;
		16'b0101111001100111: color_data = 12'b001110100111;
		16'b0101111001101000: color_data = 12'b001110100111;
		16'b0101111001110101: color_data = 12'b001110100111;
		16'b0101111001110110: color_data = 12'b001110100111;
		16'b0101111001110111: color_data = 12'b001110100111;
		16'b0101111001111000: color_data = 12'b001110100111;
		16'b0101111001111001: color_data = 12'b001110100111;
		16'b0101111001111010: color_data = 12'b001110100111;
		16'b0101111001111011: color_data = 12'b001110100111;
		16'b0101111001111100: color_data = 12'b001110100111;
		16'b0101111001111101: color_data = 12'b001110100111;
		16'b0101111001111110: color_data = 12'b001110100111;
		16'b0101111001111111: color_data = 12'b001110100111;
		16'b0101111010000000: color_data = 12'b001110100111;
		16'b0101111010001101: color_data = 12'b001110100111;
		16'b0101111010001110: color_data = 12'b001110100111;
		16'b0101111010001111: color_data = 12'b001110100111;
		16'b0101111010010000: color_data = 12'b001110100111;
		16'b0101111010010001: color_data = 12'b001110100111;
		16'b0101111010010010: color_data = 12'b001110100111;
		16'b0101111010010011: color_data = 12'b001110100111;
		16'b0101111010010100: color_data = 12'b001110100111;
		16'b0101111010010101: color_data = 12'b001110100111;
		16'b0101111010010110: color_data = 12'b001110100111;
		16'b0101111010010111: color_data = 12'b001110100111;
		16'b0101111010011000: color_data = 12'b001110100111;
		16'b0101111010011001: color_data = 12'b001110100111;
		16'b0101111010100000: color_data = 12'b001110100111;
		16'b0101111010100001: color_data = 12'b001110100111;
		16'b0101111010100010: color_data = 12'b001110100111;
		16'b0101111010100011: color_data = 12'b001110100111;
		16'b0101111010100100: color_data = 12'b001110100111;
		16'b0101111010100101: color_data = 12'b001110100111;
		16'b0101111010100110: color_data = 12'b001110100111;
		16'b0101111010100111: color_data = 12'b001110100111;
		16'b0101111010101000: color_data = 12'b001110100111;
		16'b0101111010101001: color_data = 12'b001110100111;
		16'b0101111010101010: color_data = 12'b001110100111;
		16'b0101111010101011: color_data = 12'b001110100111;
		16'b0101111011001011: color_data = 12'b001110100111;
		16'b0101111011001100: color_data = 12'b001110100111;
		16'b0101111011001101: color_data = 12'b001110100111;
		16'b0101111011001110: color_data = 12'b001110100111;
		16'b0101111011001111: color_data = 12'b001110100111;
		16'b0101111011010000: color_data = 12'b001110100111;
		16'b0101111011010001: color_data = 12'b001110100111;
		16'b0101111011010010: color_data = 12'b001110100111;
		16'b0101111011010011: color_data = 12'b001110100111;
		16'b0101111011010100: color_data = 12'b001110100111;
		16'b0101111011010101: color_data = 12'b001110100111;
		16'b0101111011010110: color_data = 12'b001110100111;
		16'b0101111011010111: color_data = 12'b001110100111;
		16'b0101111011011000: color_data = 12'b001110100111;
		16'b0101111011011001: color_data = 12'b001110100111;
		16'b0101111011011010: color_data = 12'b001110100111;
		16'b0101111011011011: color_data = 12'b001110100111;
		16'b0101111011011100: color_data = 12'b001110100111;
		16'b0101111011011101: color_data = 12'b001110100111;
		16'b0101111011011110: color_data = 12'b001110100111;
		16'b0101111011011111: color_data = 12'b001110100111;
		16'b0101111011100000: color_data = 12'b001110100111;
		16'b0101111011100001: color_data = 12'b001110100111;
		16'b0101111011100010: color_data = 12'b001110100111;
		16'b0101111011100011: color_data = 12'b001110100111;
		16'b0101111011100100: color_data = 12'b001110100111;
		16'b0101111011100101: color_data = 12'b001110100111;
		16'b0101111011100110: color_data = 12'b001110100111;
		16'b0101111011100111: color_data = 12'b001110100111;
		16'b0101111011101000: color_data = 12'b001110100111;
		16'b0101111011110110: color_data = 12'b001110100111;
		16'b0101111011110111: color_data = 12'b001110100111;
		16'b0101111011111000: color_data = 12'b001110100111;
		16'b0101111011111001: color_data = 12'b001110100111;
		16'b0101111011111010: color_data = 12'b001110100111;
		16'b0101111011111011: color_data = 12'b001110100111;
		16'b0101111011111100: color_data = 12'b001110100111;
		16'b0101111011111101: color_data = 12'b001110100111;
		16'b0101111011111110: color_data = 12'b001110100111;
		16'b0101111011111111: color_data = 12'b001110100111;
		16'b0101111100000000: color_data = 12'b001110100111;
		16'b0101111100000001: color_data = 12'b001110100111;
		16'b0101111100011010: color_data = 12'b001110100111;
		16'b0101111100011011: color_data = 12'b001110100111;
		16'b0101111100011100: color_data = 12'b001110100111;
		16'b0101111100011101: color_data = 12'b001110100111;
		16'b0101111100011110: color_data = 12'b001110100111;
		16'b0101111100011111: color_data = 12'b001110100111;
		16'b0101111100100000: color_data = 12'b001110100111;
		16'b0101111100100001: color_data = 12'b001110100111;
		16'b0101111100100010: color_data = 12'b001110100111;
		16'b0101111100100011: color_data = 12'b001110100111;
		16'b0101111100100100: color_data = 12'b001110100111;
		16'b0101111100100101: color_data = 12'b001110100111;
		16'b0101111100100110: color_data = 12'b001110100111;
		16'b0101111100101101: color_data = 12'b001110100111;
		16'b0101111100101110: color_data = 12'b001110100111;
		16'b0101111100101111: color_data = 12'b001110100111;
		16'b0101111100110000: color_data = 12'b001110100111;
		16'b0101111100110001: color_data = 12'b001110100111;
		16'b0101111100110010: color_data = 12'b001110100111;
		16'b0101111100110011: color_data = 12'b001110100111;
		16'b0101111100110100: color_data = 12'b001110100111;
		16'b0101111100110101: color_data = 12'b001110100111;
		16'b0101111100110110: color_data = 12'b001110100111;
		16'b0101111100110111: color_data = 12'b001110100111;
		16'b0101111100111000: color_data = 12'b001110100111;
		16'b0101111101000101: color_data = 12'b001110100111;
		16'b0101111101000110: color_data = 12'b001110100111;
		16'b0101111101000111: color_data = 12'b001110100111;
		16'b0101111101001000: color_data = 12'b001110100111;
		16'b0101111101001001: color_data = 12'b001110100111;
		16'b0101111101001010: color_data = 12'b001110100111;
		16'b0101111101001011: color_data = 12'b001110100111;
		16'b0101111101001100: color_data = 12'b001110100111;
		16'b0101111101001101: color_data = 12'b001110100111;
		16'b0101111101001110: color_data = 12'b001110100111;
		16'b0101111101001111: color_data = 12'b001110100111;
		16'b0101111101010000: color_data = 12'b001110100111;
		16'b0101111101010001: color_data = 12'b001110100111;
		16'b0101111101011000: color_data = 12'b001110100111;
		16'b0101111101011001: color_data = 12'b001110100111;
		16'b0101111101011010: color_data = 12'b001110100111;
		16'b0101111101011011: color_data = 12'b001110100111;
		16'b0101111101011100: color_data = 12'b001110100111;
		16'b0101111101011101: color_data = 12'b001110100111;
		16'b0101111101011110: color_data = 12'b001110100111;
		16'b0101111101011111: color_data = 12'b001110100111;
		16'b0101111101100000: color_data = 12'b001110100111;
		16'b0101111101100001: color_data = 12'b001110100111;
		16'b0101111101100010: color_data = 12'b001110100111;
		16'b0101111101100011: color_data = 12'b001110100111;
		16'b0110000000000000: color_data = 12'b001110100111;
		16'b0110000000000001: color_data = 12'b001110100111;
		16'b0110000000000010: color_data = 12'b001110100111;
		16'b0110000000000011: color_data = 12'b001110100111;
		16'b0110000000000100: color_data = 12'b001110100111;
		16'b0110000000000101: color_data = 12'b001110100111;
		16'b0110000000000110: color_data = 12'b001110100111;
		16'b0110000000000111: color_data = 12'b001110100111;
		16'b0110000000001000: color_data = 12'b001110100111;
		16'b0110000000001001: color_data = 12'b001110100111;
		16'b0110000000001010: color_data = 12'b001110100111;
		16'b0110000000001011: color_data = 12'b001110100111;
		16'b0110000000001100: color_data = 12'b001110100111;
		16'b0110000000101011: color_data = 12'b001110100111;
		16'b0110000000101100: color_data = 12'b001110100111;
		16'b0110000000101101: color_data = 12'b001110100111;
		16'b0110000000101110: color_data = 12'b001110100111;
		16'b0110000000101111: color_data = 12'b001110100111;
		16'b0110000000110000: color_data = 12'b001110100111;
		16'b0110000000110001: color_data = 12'b001110100111;
		16'b0110000000110010: color_data = 12'b001110100111;
		16'b0110000000110011: color_data = 12'b001110100111;
		16'b0110000000110100: color_data = 12'b001110100111;
		16'b0110000000110101: color_data = 12'b001110100111;
		16'b0110000000110110: color_data = 12'b001110100111;
		16'b0110000000110111: color_data = 12'b001110100111;
		16'b0110000000111000: color_data = 12'b001110100111;
		16'b0110000000111001: color_data = 12'b001110100111;
		16'b0110000000111010: color_data = 12'b001110100111;
		16'b0110000000111011: color_data = 12'b001110100111;
		16'b0110000000111100: color_data = 12'b001110100111;
		16'b0110000000111101: color_data = 12'b001110100111;
		16'b0110000000111110: color_data = 12'b001110100111;
		16'b0110000000111111: color_data = 12'b001110100111;
		16'b0110000001000000: color_data = 12'b001110100111;
		16'b0110000001000001: color_data = 12'b001110100111;
		16'b0110000001000010: color_data = 12'b001110100111;
		16'b0110000001000011: color_data = 12'b001110100111;
		16'b0110000001000100: color_data = 12'b001110100111;
		16'b0110000001000101: color_data = 12'b001110100111;
		16'b0110000001000110: color_data = 12'b001110100111;
		16'b0110000001000111: color_data = 12'b001110100111;
		16'b0110000001001000: color_data = 12'b001110100111;
		16'b0110000001001001: color_data = 12'b001110100111;
		16'b0110000001001010: color_data = 12'b001110100111;
		16'b0110000001001011: color_data = 12'b001110100111;
		16'b0110000001001100: color_data = 12'b001110100111;
		16'b0110000001001101: color_data = 12'b001110100111;
		16'b0110000001001110: color_data = 12'b001110100111;
		16'b0110000001001111: color_data = 12'b001110100111;
		16'b0110000001011100: color_data = 12'b001110100111;
		16'b0110000001011101: color_data = 12'b001110100111;
		16'b0110000001011110: color_data = 12'b001110100111;
		16'b0110000001011111: color_data = 12'b001110100111;
		16'b0110000001100000: color_data = 12'b001110100111;
		16'b0110000001100001: color_data = 12'b001110100111;
		16'b0110000001100010: color_data = 12'b001110100111;
		16'b0110000001100011: color_data = 12'b001110100111;
		16'b0110000001100100: color_data = 12'b001110100111;
		16'b0110000001100101: color_data = 12'b001110100111;
		16'b0110000001100110: color_data = 12'b001110100111;
		16'b0110000001100111: color_data = 12'b001110100111;
		16'b0110000001101000: color_data = 12'b001110100111;
		16'b0110000001110101: color_data = 12'b001110100111;
		16'b0110000001110110: color_data = 12'b001110100111;
		16'b0110000001110111: color_data = 12'b001110100111;
		16'b0110000001111000: color_data = 12'b001110100111;
		16'b0110000001111001: color_data = 12'b001110100111;
		16'b0110000001111010: color_data = 12'b001110100111;
		16'b0110000001111011: color_data = 12'b001110100111;
		16'b0110000001111100: color_data = 12'b001110100111;
		16'b0110000001111101: color_data = 12'b001110100111;
		16'b0110000001111110: color_data = 12'b001110100111;
		16'b0110000001111111: color_data = 12'b001110100111;
		16'b0110000010000000: color_data = 12'b001110100111;
		16'b0110000010001101: color_data = 12'b001110100111;
		16'b0110000010001110: color_data = 12'b001110100111;
		16'b0110000010001111: color_data = 12'b001110100111;
		16'b0110000010010000: color_data = 12'b001110100111;
		16'b0110000010010001: color_data = 12'b001110100111;
		16'b0110000010010010: color_data = 12'b001110100111;
		16'b0110000010010011: color_data = 12'b001110100111;
		16'b0110000010010100: color_data = 12'b001110100111;
		16'b0110000010010101: color_data = 12'b001110100111;
		16'b0110000010010110: color_data = 12'b001110100111;
		16'b0110000010010111: color_data = 12'b001110100111;
		16'b0110000010011000: color_data = 12'b001110100111;
		16'b0110000010011001: color_data = 12'b001110100111;
		16'b0110000010100000: color_data = 12'b001110100111;
		16'b0110000010100001: color_data = 12'b001110100111;
		16'b0110000010100010: color_data = 12'b001110100111;
		16'b0110000010100011: color_data = 12'b001110100111;
		16'b0110000010100100: color_data = 12'b001110100111;
		16'b0110000010100101: color_data = 12'b001110100111;
		16'b0110000010100110: color_data = 12'b001110100111;
		16'b0110000010100111: color_data = 12'b001110100111;
		16'b0110000010101000: color_data = 12'b001110100111;
		16'b0110000010101001: color_data = 12'b001110100111;
		16'b0110000010101010: color_data = 12'b001110100111;
		16'b0110000010101011: color_data = 12'b001110100111;
		16'b0110000011001011: color_data = 12'b001110100111;
		16'b0110000011001100: color_data = 12'b001110100111;
		16'b0110000011001101: color_data = 12'b001110100111;
		16'b0110000011001110: color_data = 12'b001110100111;
		16'b0110000011001111: color_data = 12'b001110100111;
		16'b0110000011010000: color_data = 12'b001110100111;
		16'b0110000011010001: color_data = 12'b001110100111;
		16'b0110000011010010: color_data = 12'b001110100111;
		16'b0110000011010011: color_data = 12'b001110100111;
		16'b0110000011010100: color_data = 12'b001110100111;
		16'b0110000011010101: color_data = 12'b001110100111;
		16'b0110000011010110: color_data = 12'b001110100111;
		16'b0110000011010111: color_data = 12'b001110100111;
		16'b0110000011011000: color_data = 12'b001110100111;
		16'b0110000011011001: color_data = 12'b001110100111;
		16'b0110000011011010: color_data = 12'b001110100111;
		16'b0110000011011011: color_data = 12'b001110100111;
		16'b0110000011011100: color_data = 12'b001110100111;
		16'b0110000011011101: color_data = 12'b001110100111;
		16'b0110000011011110: color_data = 12'b001110100111;
		16'b0110000011011111: color_data = 12'b001110100111;
		16'b0110000011100000: color_data = 12'b001110100111;
		16'b0110000011100001: color_data = 12'b001110100111;
		16'b0110000011100010: color_data = 12'b001110100111;
		16'b0110000011100011: color_data = 12'b001110100111;
		16'b0110000011100100: color_data = 12'b001110100111;
		16'b0110000011100101: color_data = 12'b001110100111;
		16'b0110000011100110: color_data = 12'b001110100111;
		16'b0110000011100111: color_data = 12'b001110100111;
		16'b0110000011101000: color_data = 12'b001110100111;
		16'b0110000011110110: color_data = 12'b001110100111;
		16'b0110000011110111: color_data = 12'b001110100111;
		16'b0110000011111000: color_data = 12'b001110100111;
		16'b0110000011111001: color_data = 12'b001110100111;
		16'b0110000011111010: color_data = 12'b001110100111;
		16'b0110000011111011: color_data = 12'b001110100111;
		16'b0110000011111100: color_data = 12'b001110100111;
		16'b0110000011111101: color_data = 12'b001110100111;
		16'b0110000011111110: color_data = 12'b001110100111;
		16'b0110000011111111: color_data = 12'b001110100111;
		16'b0110000100000000: color_data = 12'b001110100111;
		16'b0110000100000001: color_data = 12'b001110100111;
		16'b0110000100011010: color_data = 12'b001110100111;
		16'b0110000100011011: color_data = 12'b001110100111;
		16'b0110000100011100: color_data = 12'b001110100111;
		16'b0110000100011101: color_data = 12'b001110100111;
		16'b0110000100011110: color_data = 12'b001110100111;
		16'b0110000100011111: color_data = 12'b001110100111;
		16'b0110000100100000: color_data = 12'b001110100111;
		16'b0110000100100001: color_data = 12'b001110100111;
		16'b0110000100100010: color_data = 12'b001110100111;
		16'b0110000100100011: color_data = 12'b001110100111;
		16'b0110000100100100: color_data = 12'b001110100111;
		16'b0110000100100101: color_data = 12'b001110100111;
		16'b0110000100100110: color_data = 12'b001110100111;
		16'b0110000100101101: color_data = 12'b001110100111;
		16'b0110000100101110: color_data = 12'b001110100111;
		16'b0110000100101111: color_data = 12'b001110100111;
		16'b0110000100110000: color_data = 12'b001110100111;
		16'b0110000100110001: color_data = 12'b001110100111;
		16'b0110000100110010: color_data = 12'b001110100111;
		16'b0110000100110011: color_data = 12'b001110100111;
		16'b0110000100110100: color_data = 12'b001110100111;
		16'b0110000100110101: color_data = 12'b001110100111;
		16'b0110000100110110: color_data = 12'b001110100111;
		16'b0110000100110111: color_data = 12'b001110100111;
		16'b0110000100111000: color_data = 12'b001110100111;
		16'b0110000101000101: color_data = 12'b001110100111;
		16'b0110000101000110: color_data = 12'b001110100111;
		16'b0110000101000111: color_data = 12'b001110100111;
		16'b0110000101001000: color_data = 12'b001110100111;
		16'b0110000101001001: color_data = 12'b001110100111;
		16'b0110000101001010: color_data = 12'b001110100111;
		16'b0110000101001011: color_data = 12'b001110100111;
		16'b0110000101001100: color_data = 12'b001110100111;
		16'b0110000101001101: color_data = 12'b001110100111;
		16'b0110000101001110: color_data = 12'b001110100111;
		16'b0110000101001111: color_data = 12'b001110100111;
		16'b0110000101010000: color_data = 12'b001110100111;
		16'b0110000101010001: color_data = 12'b001110100111;
		16'b0110000101011000: color_data = 12'b001110100111;
		16'b0110000101011001: color_data = 12'b001110100111;
		16'b0110000101011010: color_data = 12'b001110100111;
		16'b0110000101011011: color_data = 12'b001110100111;
		16'b0110000101011100: color_data = 12'b001110100111;
		16'b0110000101011101: color_data = 12'b001110100111;
		16'b0110000101011110: color_data = 12'b001110100111;
		16'b0110000101011111: color_data = 12'b001110100111;
		16'b0110000101100000: color_data = 12'b001110100111;
		16'b0110000101100001: color_data = 12'b001110100111;
		16'b0110000101100010: color_data = 12'b001110100111;
		16'b0110000101100011: color_data = 12'b001110100111;
		16'b0110001000000000: color_data = 12'b001110100111;
		16'b0110001000000001: color_data = 12'b001110100111;
		16'b0110001000000010: color_data = 12'b001110100111;
		16'b0110001000000011: color_data = 12'b001110100111;
		16'b0110001000000100: color_data = 12'b001110100111;
		16'b0110001000000101: color_data = 12'b001110100111;
		16'b0110001000000110: color_data = 12'b001110100111;
		16'b0110001000000111: color_data = 12'b001110100111;
		16'b0110001000001000: color_data = 12'b001110100111;
		16'b0110001000001001: color_data = 12'b001110100111;
		16'b0110001000001010: color_data = 12'b001110100111;
		16'b0110001000001011: color_data = 12'b001110100111;
		16'b0110001000001100: color_data = 12'b001110100111;
		16'b0110001000101011: color_data = 12'b001110100111;
		16'b0110001000101100: color_data = 12'b001110100111;
		16'b0110001000101101: color_data = 12'b001110100111;
		16'b0110001000101110: color_data = 12'b001110100111;
		16'b0110001000101111: color_data = 12'b001110100111;
		16'b0110001000110000: color_data = 12'b001110100111;
		16'b0110001000110001: color_data = 12'b001110100111;
		16'b0110001000110010: color_data = 12'b001110100111;
		16'b0110001000110011: color_data = 12'b001110100111;
		16'b0110001000110100: color_data = 12'b001110100111;
		16'b0110001000110101: color_data = 12'b001110100111;
		16'b0110001000110110: color_data = 12'b001110100111;
		16'b0110001000110111: color_data = 12'b001110100111;
		16'b0110001000111000: color_data = 12'b001110100111;
		16'b0110001000111001: color_data = 12'b001110100111;
		16'b0110001000111010: color_data = 12'b001110100111;
		16'b0110001000111011: color_data = 12'b001110100111;
		16'b0110001000111100: color_data = 12'b001110100111;
		16'b0110001000111101: color_data = 12'b001110100111;
		16'b0110001000111110: color_data = 12'b001110100111;
		16'b0110001000111111: color_data = 12'b001110100111;
		16'b0110001001000000: color_data = 12'b001110100111;
		16'b0110001001000001: color_data = 12'b001110100111;
		16'b0110001001000010: color_data = 12'b001110100111;
		16'b0110001001000011: color_data = 12'b001110100111;
		16'b0110001001000100: color_data = 12'b001110100111;
		16'b0110001001000101: color_data = 12'b001110100111;
		16'b0110001001000110: color_data = 12'b001110100111;
		16'b0110001001000111: color_data = 12'b001110100111;
		16'b0110001001001000: color_data = 12'b001110100111;
		16'b0110001001001001: color_data = 12'b001110100111;
		16'b0110001001001010: color_data = 12'b001110100111;
		16'b0110001001001011: color_data = 12'b001110100111;
		16'b0110001001001100: color_data = 12'b001110100111;
		16'b0110001001001101: color_data = 12'b001110100111;
		16'b0110001001001110: color_data = 12'b001110100111;
		16'b0110001001001111: color_data = 12'b001110100111;
		16'b0110001001011100: color_data = 12'b001110100111;
		16'b0110001001011101: color_data = 12'b001110100111;
		16'b0110001001011110: color_data = 12'b001110100111;
		16'b0110001001011111: color_data = 12'b001110100111;
		16'b0110001001100000: color_data = 12'b001110100111;
		16'b0110001001100001: color_data = 12'b001110100111;
		16'b0110001001100010: color_data = 12'b001110100111;
		16'b0110001001100011: color_data = 12'b001110100111;
		16'b0110001001100100: color_data = 12'b001110100111;
		16'b0110001001100101: color_data = 12'b001110100111;
		16'b0110001001100110: color_data = 12'b001110100111;
		16'b0110001001100111: color_data = 12'b001110100111;
		16'b0110001001101000: color_data = 12'b001110100111;
		16'b0110001001110101: color_data = 12'b001110100111;
		16'b0110001001110110: color_data = 12'b001110100111;
		16'b0110001001110111: color_data = 12'b001110100111;
		16'b0110001001111000: color_data = 12'b001110100111;
		16'b0110001001111001: color_data = 12'b001110100111;
		16'b0110001001111010: color_data = 12'b001110100111;
		16'b0110001001111011: color_data = 12'b001110100111;
		16'b0110001001111100: color_data = 12'b001110100111;
		16'b0110001001111101: color_data = 12'b001110100111;
		16'b0110001001111110: color_data = 12'b001110100111;
		16'b0110001001111111: color_data = 12'b001110100111;
		16'b0110001010000000: color_data = 12'b001110100111;
		16'b0110001010001101: color_data = 12'b001110100111;
		16'b0110001010001110: color_data = 12'b001110100111;
		16'b0110001010001111: color_data = 12'b001110100111;
		16'b0110001010010000: color_data = 12'b001110100111;
		16'b0110001010010001: color_data = 12'b001110100111;
		16'b0110001010010010: color_data = 12'b001110100111;
		16'b0110001010010011: color_data = 12'b001110100111;
		16'b0110001010010100: color_data = 12'b001110100111;
		16'b0110001010010101: color_data = 12'b001110100111;
		16'b0110001010010110: color_data = 12'b001110100111;
		16'b0110001010010111: color_data = 12'b001110100111;
		16'b0110001010011000: color_data = 12'b001110100111;
		16'b0110001010011001: color_data = 12'b001110100111;
		16'b0110001010100000: color_data = 12'b001110100111;
		16'b0110001010100001: color_data = 12'b001110100111;
		16'b0110001010100010: color_data = 12'b001110100111;
		16'b0110001010100011: color_data = 12'b001110100111;
		16'b0110001010100100: color_data = 12'b001110100111;
		16'b0110001010100101: color_data = 12'b001110100111;
		16'b0110001010100110: color_data = 12'b001110100111;
		16'b0110001010100111: color_data = 12'b001110100111;
		16'b0110001010101000: color_data = 12'b001110100111;
		16'b0110001010101001: color_data = 12'b001110100111;
		16'b0110001010101010: color_data = 12'b001110100111;
		16'b0110001010101011: color_data = 12'b001110100111;
		16'b0110001011001011: color_data = 12'b001110100111;
		16'b0110001011001100: color_data = 12'b001110100111;
		16'b0110001011001101: color_data = 12'b001110100111;
		16'b0110001011001110: color_data = 12'b001110100111;
		16'b0110001011001111: color_data = 12'b001110100111;
		16'b0110001011010000: color_data = 12'b001110100111;
		16'b0110001011010001: color_data = 12'b001110100111;
		16'b0110001011010010: color_data = 12'b001110100111;
		16'b0110001011010011: color_data = 12'b001110100111;
		16'b0110001011010100: color_data = 12'b001110100111;
		16'b0110001011010101: color_data = 12'b001110100111;
		16'b0110001011010110: color_data = 12'b001110100111;
		16'b0110001011010111: color_data = 12'b001110100111;
		16'b0110001011011000: color_data = 12'b001110100111;
		16'b0110001011011001: color_data = 12'b001110100111;
		16'b0110001011011010: color_data = 12'b001110100111;
		16'b0110001011011011: color_data = 12'b001110100111;
		16'b0110001011011100: color_data = 12'b001110100111;
		16'b0110001011011101: color_data = 12'b001110100111;
		16'b0110001011011110: color_data = 12'b001110100111;
		16'b0110001011011111: color_data = 12'b001110100111;
		16'b0110001011100000: color_data = 12'b001110100111;
		16'b0110001011100001: color_data = 12'b001110100111;
		16'b0110001011100010: color_data = 12'b001110100111;
		16'b0110001011100011: color_data = 12'b001110100111;
		16'b0110001011100100: color_data = 12'b001110100111;
		16'b0110001011100101: color_data = 12'b001110100111;
		16'b0110001011100110: color_data = 12'b001110100111;
		16'b0110001011100111: color_data = 12'b001110100111;
		16'b0110001011101000: color_data = 12'b001110100111;
		16'b0110001011110110: color_data = 12'b001110100111;
		16'b0110001011110111: color_data = 12'b001110100111;
		16'b0110001011111000: color_data = 12'b001110100111;
		16'b0110001011111001: color_data = 12'b001110100111;
		16'b0110001011111010: color_data = 12'b001110100111;
		16'b0110001011111011: color_data = 12'b001110100111;
		16'b0110001011111100: color_data = 12'b001110100111;
		16'b0110001011111101: color_data = 12'b001110100111;
		16'b0110001011111110: color_data = 12'b001110100111;
		16'b0110001011111111: color_data = 12'b001110100111;
		16'b0110001100000000: color_data = 12'b001110100111;
		16'b0110001100000001: color_data = 12'b001110100111;
		16'b0110001100011010: color_data = 12'b001110100111;
		16'b0110001100011011: color_data = 12'b001110100111;
		16'b0110001100011100: color_data = 12'b001110100111;
		16'b0110001100011101: color_data = 12'b001110100111;
		16'b0110001100011110: color_data = 12'b001110100111;
		16'b0110001100011111: color_data = 12'b001110100111;
		16'b0110001100100000: color_data = 12'b001110100111;
		16'b0110001100100001: color_data = 12'b001110100111;
		16'b0110001100100010: color_data = 12'b001110100111;
		16'b0110001100100011: color_data = 12'b001110100111;
		16'b0110001100100100: color_data = 12'b001110100111;
		16'b0110001100100101: color_data = 12'b001110100111;
		16'b0110001100100110: color_data = 12'b001110100111;
		16'b0110001100101101: color_data = 12'b001110100111;
		16'b0110001100101110: color_data = 12'b001110100111;
		16'b0110001100101111: color_data = 12'b001110100111;
		16'b0110001100110000: color_data = 12'b001110100111;
		16'b0110001100110001: color_data = 12'b001110100111;
		16'b0110001100110010: color_data = 12'b001110100111;
		16'b0110001100110011: color_data = 12'b001110100111;
		16'b0110001100110100: color_data = 12'b001110100111;
		16'b0110001100110101: color_data = 12'b001110100111;
		16'b0110001100110110: color_data = 12'b001110100111;
		16'b0110001100110111: color_data = 12'b001110100111;
		16'b0110001100111000: color_data = 12'b001110100111;
		16'b0110001101000101: color_data = 12'b001110100111;
		16'b0110001101000110: color_data = 12'b001110100111;
		16'b0110001101000111: color_data = 12'b001110100111;
		16'b0110001101001000: color_data = 12'b001110100111;
		16'b0110001101001001: color_data = 12'b001110100111;
		16'b0110001101001010: color_data = 12'b001110100111;
		16'b0110001101001011: color_data = 12'b001110100111;
		16'b0110001101001100: color_data = 12'b001110100111;
		16'b0110001101001101: color_data = 12'b001110100111;
		16'b0110001101001110: color_data = 12'b001110100111;
		16'b0110001101001111: color_data = 12'b001110100111;
		16'b0110001101010000: color_data = 12'b001110100111;
		16'b0110001101010001: color_data = 12'b001110100111;
		16'b0110001101011000: color_data = 12'b001110100111;
		16'b0110001101011001: color_data = 12'b001110100111;
		16'b0110001101011010: color_data = 12'b001110100111;
		16'b0110001101011011: color_data = 12'b001110100111;
		16'b0110001101011100: color_data = 12'b001110100111;
		16'b0110001101011101: color_data = 12'b001110100111;
		16'b0110001101011110: color_data = 12'b001110100111;
		16'b0110001101011111: color_data = 12'b001110100111;
		16'b0110001101100000: color_data = 12'b001110100111;
		16'b0110001101100001: color_data = 12'b001110100111;
		16'b0110001101100010: color_data = 12'b001110100111;
		16'b0110001101100011: color_data = 12'b001110100111;
		16'b0110010000000000: color_data = 12'b001110100111;
		16'b0110010000000001: color_data = 12'b001110100111;
		16'b0110010000000010: color_data = 12'b001110100111;
		16'b0110010000000011: color_data = 12'b001110100111;
		16'b0110010000000100: color_data = 12'b001110100111;
		16'b0110010000000101: color_data = 12'b001110100111;
		16'b0110010000000110: color_data = 12'b001110100111;
		16'b0110010000000111: color_data = 12'b001110100111;
		16'b0110010000001000: color_data = 12'b001110100111;
		16'b0110010000001001: color_data = 12'b001110100111;
		16'b0110010000001010: color_data = 12'b001110100111;
		16'b0110010000001011: color_data = 12'b001110100111;
		16'b0110010000001100: color_data = 12'b001110100111;
		16'b0110010000101011: color_data = 12'b001110100111;
		16'b0110010000101100: color_data = 12'b001110100111;
		16'b0110010000101101: color_data = 12'b001110100111;
		16'b0110010000101110: color_data = 12'b001110100111;
		16'b0110010000101111: color_data = 12'b001110100111;
		16'b0110010000110000: color_data = 12'b001110100111;
		16'b0110010000110001: color_data = 12'b001110100111;
		16'b0110010000110010: color_data = 12'b001110100111;
		16'b0110010000110011: color_data = 12'b001110100111;
		16'b0110010000110100: color_data = 12'b001110100111;
		16'b0110010000110101: color_data = 12'b001110100111;
		16'b0110010000110110: color_data = 12'b001110100111;
		16'b0110010000110111: color_data = 12'b001110100111;
		16'b0110010000111000: color_data = 12'b001110100111;
		16'b0110010000111001: color_data = 12'b001110100111;
		16'b0110010000111010: color_data = 12'b001110100111;
		16'b0110010000111011: color_data = 12'b001110100111;
		16'b0110010000111100: color_data = 12'b001110100111;
		16'b0110010000111101: color_data = 12'b001110100111;
		16'b0110010000111110: color_data = 12'b001110100111;
		16'b0110010000111111: color_data = 12'b001110100111;
		16'b0110010001000000: color_data = 12'b001110100111;
		16'b0110010001000001: color_data = 12'b001110100111;
		16'b0110010001000010: color_data = 12'b001110100111;
		16'b0110010001000011: color_data = 12'b001110100111;
		16'b0110010001000100: color_data = 12'b001110100111;
		16'b0110010001000101: color_data = 12'b001110100111;
		16'b0110010001000110: color_data = 12'b001110100111;
		16'b0110010001000111: color_data = 12'b001110100111;
		16'b0110010001001000: color_data = 12'b001110100111;
		16'b0110010001001001: color_data = 12'b001110100111;
		16'b0110010001001010: color_data = 12'b001110100111;
		16'b0110010001001011: color_data = 12'b001110100111;
		16'b0110010001001100: color_data = 12'b001110100111;
		16'b0110010001001101: color_data = 12'b001110100111;
		16'b0110010001001110: color_data = 12'b001110100111;
		16'b0110010001001111: color_data = 12'b001110100111;
		16'b0110010001011100: color_data = 12'b001110100111;
		16'b0110010001011101: color_data = 12'b001110100111;
		16'b0110010001011110: color_data = 12'b001110100111;
		16'b0110010001011111: color_data = 12'b001110100111;
		16'b0110010001100000: color_data = 12'b001110100111;
		16'b0110010001100001: color_data = 12'b001110100111;
		16'b0110010001100010: color_data = 12'b001110100111;
		16'b0110010001100011: color_data = 12'b001110100111;
		16'b0110010001100100: color_data = 12'b001110100111;
		16'b0110010001100101: color_data = 12'b001110100111;
		16'b0110010001100110: color_data = 12'b001110100111;
		16'b0110010001100111: color_data = 12'b001110100111;
		16'b0110010001101000: color_data = 12'b001110100111;
		16'b0110010001110101: color_data = 12'b001110100111;
		16'b0110010001110110: color_data = 12'b001110100111;
		16'b0110010001110111: color_data = 12'b001110100111;
		16'b0110010001111000: color_data = 12'b001110100111;
		16'b0110010001111001: color_data = 12'b001110100111;
		16'b0110010001111010: color_data = 12'b001110100111;
		16'b0110010001111011: color_data = 12'b001110100111;
		16'b0110010001111100: color_data = 12'b001110100111;
		16'b0110010001111101: color_data = 12'b001110100111;
		16'b0110010001111110: color_data = 12'b001110100111;
		16'b0110010001111111: color_data = 12'b001110100111;
		16'b0110010010000000: color_data = 12'b001110100111;
		16'b0110010010001101: color_data = 12'b001110100111;
		16'b0110010010001110: color_data = 12'b001110100111;
		16'b0110010010001111: color_data = 12'b001110100111;
		16'b0110010010010000: color_data = 12'b001110100111;
		16'b0110010010010001: color_data = 12'b001110100111;
		16'b0110010010010010: color_data = 12'b001110100111;
		16'b0110010010010011: color_data = 12'b001110100111;
		16'b0110010010010100: color_data = 12'b001110100111;
		16'b0110010010010101: color_data = 12'b001110100111;
		16'b0110010010010110: color_data = 12'b001110100111;
		16'b0110010010010111: color_data = 12'b001110100111;
		16'b0110010010011000: color_data = 12'b001110100111;
		16'b0110010010011001: color_data = 12'b001110100111;
		16'b0110010010100000: color_data = 12'b001110100111;
		16'b0110010010100001: color_data = 12'b001110100111;
		16'b0110010010100010: color_data = 12'b001110100111;
		16'b0110010010100011: color_data = 12'b001110100111;
		16'b0110010010100100: color_data = 12'b001110100111;
		16'b0110010010100101: color_data = 12'b001110100111;
		16'b0110010010100110: color_data = 12'b001110100111;
		16'b0110010010100111: color_data = 12'b001110100111;
		16'b0110010010101000: color_data = 12'b001110100111;
		16'b0110010010101001: color_data = 12'b001110100111;
		16'b0110010010101010: color_data = 12'b001110100111;
		16'b0110010010101011: color_data = 12'b001110100111;
		16'b0110010011001011: color_data = 12'b001110100111;
		16'b0110010011001100: color_data = 12'b001110100111;
		16'b0110010011001101: color_data = 12'b001110100111;
		16'b0110010011001110: color_data = 12'b001110100111;
		16'b0110010011001111: color_data = 12'b001110100111;
		16'b0110010011010000: color_data = 12'b001110100111;
		16'b0110010011010001: color_data = 12'b001110100111;
		16'b0110010011010010: color_data = 12'b001110100111;
		16'b0110010011010011: color_data = 12'b001110100111;
		16'b0110010011010100: color_data = 12'b001110100111;
		16'b0110010011010101: color_data = 12'b001110100111;
		16'b0110010011010110: color_data = 12'b001110100111;
		16'b0110010011010111: color_data = 12'b001110100111;
		16'b0110010011011000: color_data = 12'b001110100111;
		16'b0110010011011001: color_data = 12'b001110100111;
		16'b0110010011011010: color_data = 12'b001110100111;
		16'b0110010011011011: color_data = 12'b001110100111;
		16'b0110010011011100: color_data = 12'b001110100111;
		16'b0110010011011101: color_data = 12'b001110100111;
		16'b0110010011011110: color_data = 12'b001110100111;
		16'b0110010011011111: color_data = 12'b001110100111;
		16'b0110010011100000: color_data = 12'b001110100111;
		16'b0110010011100001: color_data = 12'b001110100111;
		16'b0110010011100010: color_data = 12'b001110100111;
		16'b0110010011100011: color_data = 12'b001110100111;
		16'b0110010011100100: color_data = 12'b001110100111;
		16'b0110010011100101: color_data = 12'b001110100111;
		16'b0110010011100110: color_data = 12'b001110100111;
		16'b0110010011100111: color_data = 12'b001110100111;
		16'b0110010011101000: color_data = 12'b001110100111;
		16'b0110010011110110: color_data = 12'b001110100111;
		16'b0110010011110111: color_data = 12'b001110100111;
		16'b0110010011111000: color_data = 12'b001110100111;
		16'b0110010011111001: color_data = 12'b001110100111;
		16'b0110010011111010: color_data = 12'b001110100111;
		16'b0110010011111011: color_data = 12'b001110100111;
		16'b0110010011111100: color_data = 12'b001110100111;
		16'b0110010011111101: color_data = 12'b001110100111;
		16'b0110010011111110: color_data = 12'b001110100111;
		16'b0110010011111111: color_data = 12'b001110100111;
		16'b0110010100000000: color_data = 12'b001110100111;
		16'b0110010100000001: color_data = 12'b001110100111;
		16'b0110010100011010: color_data = 12'b001110100111;
		16'b0110010100011011: color_data = 12'b001110100111;
		16'b0110010100011100: color_data = 12'b001110100111;
		16'b0110010100011101: color_data = 12'b001110100111;
		16'b0110010100011110: color_data = 12'b001110100111;
		16'b0110010100011111: color_data = 12'b001110100111;
		16'b0110010100100000: color_data = 12'b001110100111;
		16'b0110010100100001: color_data = 12'b001110100111;
		16'b0110010100100010: color_data = 12'b001110100111;
		16'b0110010100100011: color_data = 12'b001110100111;
		16'b0110010100100100: color_data = 12'b001110100111;
		16'b0110010100100101: color_data = 12'b001110100111;
		16'b0110010100100110: color_data = 12'b001110100111;
		16'b0110010100101101: color_data = 12'b001110100111;
		16'b0110010100101110: color_data = 12'b001110100111;
		16'b0110010100101111: color_data = 12'b001110100111;
		16'b0110010100110000: color_data = 12'b001110100111;
		16'b0110010100110001: color_data = 12'b001110100111;
		16'b0110010100110010: color_data = 12'b001110100111;
		16'b0110010100110011: color_data = 12'b001110100111;
		16'b0110010100110100: color_data = 12'b001110100111;
		16'b0110010100110101: color_data = 12'b001110100111;
		16'b0110010100110110: color_data = 12'b001110100111;
		16'b0110010100110111: color_data = 12'b001110100111;
		16'b0110010100111000: color_data = 12'b001110100111;
		16'b0110010101000101: color_data = 12'b001110100111;
		16'b0110010101000110: color_data = 12'b001110100111;
		16'b0110010101000111: color_data = 12'b001110100111;
		16'b0110010101001000: color_data = 12'b001110100111;
		16'b0110010101001001: color_data = 12'b001110100111;
		16'b0110010101001010: color_data = 12'b001110100111;
		16'b0110010101001011: color_data = 12'b001110100111;
		16'b0110010101001100: color_data = 12'b001110100111;
		16'b0110010101001101: color_data = 12'b001110100111;
		16'b0110010101001110: color_data = 12'b001110100111;
		16'b0110010101001111: color_data = 12'b001110100111;
		16'b0110010101010000: color_data = 12'b001110100111;
		16'b0110010101010001: color_data = 12'b001110100111;
		16'b0110010101011000: color_data = 12'b001110100111;
		16'b0110010101011001: color_data = 12'b001110100111;
		16'b0110010101011010: color_data = 12'b001110100111;
		16'b0110010101011011: color_data = 12'b001110100111;
		16'b0110010101011100: color_data = 12'b001110100111;
		16'b0110010101011101: color_data = 12'b001110100111;
		16'b0110010101011110: color_data = 12'b001110100111;
		16'b0110010101011111: color_data = 12'b001110100111;
		16'b0110010101100000: color_data = 12'b001110100111;
		16'b0110010101100001: color_data = 12'b001110100111;
		16'b0110010101100010: color_data = 12'b001110100111;
		16'b0110010101100011: color_data = 12'b001110100111;
		16'b0110011000000000: color_data = 12'b001110100111;
		16'b0110011000000001: color_data = 12'b001110100111;
		16'b0110011000000010: color_data = 12'b001110100111;
		16'b0110011000000011: color_data = 12'b001110100111;
		16'b0110011000000100: color_data = 12'b001110100111;
		16'b0110011000000101: color_data = 12'b001110100111;
		16'b0110011000000110: color_data = 12'b001110100111;
		16'b0110011000000111: color_data = 12'b001110100111;
		16'b0110011000001000: color_data = 12'b001110100111;
		16'b0110011000001001: color_data = 12'b001110100111;
		16'b0110011000001010: color_data = 12'b001110100111;
		16'b0110011000001011: color_data = 12'b001110100111;
		16'b0110011000001100: color_data = 12'b001110100111;
		16'b0110011000101011: color_data = 12'b001110100111;
		16'b0110011000101100: color_data = 12'b001110100111;
		16'b0110011000101101: color_data = 12'b001110100111;
		16'b0110011000101110: color_data = 12'b001110100111;
		16'b0110011000101111: color_data = 12'b001110100111;
		16'b0110011000110000: color_data = 12'b001110100111;
		16'b0110011000110001: color_data = 12'b001110100111;
		16'b0110011000110010: color_data = 12'b001110100111;
		16'b0110011000110011: color_data = 12'b001110100111;
		16'b0110011000110100: color_data = 12'b001110100111;
		16'b0110011000110101: color_data = 12'b001110100111;
		16'b0110011000110110: color_data = 12'b001110100111;
		16'b0110011000110111: color_data = 12'b001110100111;
		16'b0110011000111000: color_data = 12'b001110100111;
		16'b0110011000111001: color_data = 12'b001110100111;
		16'b0110011000111010: color_data = 12'b001110100111;
		16'b0110011000111011: color_data = 12'b001110100111;
		16'b0110011000111100: color_data = 12'b001110100111;
		16'b0110011000111101: color_data = 12'b001110100111;
		16'b0110011000111110: color_data = 12'b001110100111;
		16'b0110011000111111: color_data = 12'b001110100111;
		16'b0110011001000000: color_data = 12'b001110100111;
		16'b0110011001000001: color_data = 12'b001110100111;
		16'b0110011001000010: color_data = 12'b001110100111;
		16'b0110011001000011: color_data = 12'b001110100111;
		16'b0110011001000100: color_data = 12'b001110100111;
		16'b0110011001000101: color_data = 12'b001110100111;
		16'b0110011001000110: color_data = 12'b001110100111;
		16'b0110011001000111: color_data = 12'b001110100111;
		16'b0110011001001000: color_data = 12'b001110100111;
		16'b0110011001001001: color_data = 12'b001110100111;
		16'b0110011001001010: color_data = 12'b001110100111;
		16'b0110011001001011: color_data = 12'b001110100111;
		16'b0110011001001100: color_data = 12'b001110100111;
		16'b0110011001001101: color_data = 12'b001110100111;
		16'b0110011001001110: color_data = 12'b001110100111;
		16'b0110011001001111: color_data = 12'b001110100111;
		16'b0110011001011100: color_data = 12'b001110100111;
		16'b0110011001011101: color_data = 12'b001110100111;
		16'b0110011001011110: color_data = 12'b001110100111;
		16'b0110011001011111: color_data = 12'b001110100111;
		16'b0110011001100000: color_data = 12'b001110100111;
		16'b0110011001100001: color_data = 12'b001110100111;
		16'b0110011001100010: color_data = 12'b001110100111;
		16'b0110011001100011: color_data = 12'b001110100111;
		16'b0110011001100100: color_data = 12'b001110100111;
		16'b0110011001100101: color_data = 12'b001110100111;
		16'b0110011001100110: color_data = 12'b001110100111;
		16'b0110011001100111: color_data = 12'b001110100111;
		16'b0110011001101000: color_data = 12'b001110100111;
		16'b0110011001110101: color_data = 12'b001110100111;
		16'b0110011001110110: color_data = 12'b001110100111;
		16'b0110011001110111: color_data = 12'b001110100111;
		16'b0110011001111000: color_data = 12'b001110100111;
		16'b0110011001111001: color_data = 12'b001110100111;
		16'b0110011001111010: color_data = 12'b001110100111;
		16'b0110011001111011: color_data = 12'b001110100111;
		16'b0110011001111100: color_data = 12'b001110100111;
		16'b0110011001111101: color_data = 12'b001110100111;
		16'b0110011001111110: color_data = 12'b001110100111;
		16'b0110011001111111: color_data = 12'b001110100111;
		16'b0110011010000000: color_data = 12'b001110100111;
		16'b0110011010001101: color_data = 12'b001110100111;
		16'b0110011010001110: color_data = 12'b001110100111;
		16'b0110011010001111: color_data = 12'b001110100111;
		16'b0110011010010000: color_data = 12'b001110100111;
		16'b0110011010010001: color_data = 12'b001110100111;
		16'b0110011010010010: color_data = 12'b001110100111;
		16'b0110011010010011: color_data = 12'b001110100111;
		16'b0110011010010100: color_data = 12'b001110100111;
		16'b0110011010010101: color_data = 12'b001110100111;
		16'b0110011010010110: color_data = 12'b001110100111;
		16'b0110011010010111: color_data = 12'b001110100111;
		16'b0110011010011000: color_data = 12'b001110100111;
		16'b0110011010011001: color_data = 12'b001110100111;
		16'b0110011010100000: color_data = 12'b001110100111;
		16'b0110011010100001: color_data = 12'b001110100111;
		16'b0110011010100010: color_data = 12'b001110100111;
		16'b0110011010100011: color_data = 12'b001110100111;
		16'b0110011010100100: color_data = 12'b001110100111;
		16'b0110011010100101: color_data = 12'b001110100111;
		16'b0110011010100110: color_data = 12'b001110100111;
		16'b0110011010100111: color_data = 12'b001110100111;
		16'b0110011010101000: color_data = 12'b001110100111;
		16'b0110011010101001: color_data = 12'b001110100111;
		16'b0110011010101010: color_data = 12'b001110100111;
		16'b0110011010101011: color_data = 12'b001110100111;
		16'b0110011010111000: color_data = 12'b001110100111;
		16'b0110011010111001: color_data = 12'b001110100111;
		16'b0110011010111010: color_data = 12'b001110100111;
		16'b0110011010111011: color_data = 12'b001110100111;
		16'b0110011010111100: color_data = 12'b001110100111;
		16'b0110011010111101: color_data = 12'b001110100111;
		16'b0110011010111110: color_data = 12'b001110100111;
		16'b0110011010111111: color_data = 12'b001110100111;
		16'b0110011011000000: color_data = 12'b001110100111;
		16'b0110011011000001: color_data = 12'b001110100111;
		16'b0110011011000010: color_data = 12'b001110100111;
		16'b0110011011000011: color_data = 12'b001110100111;
		16'b0110011011000100: color_data = 12'b001110100111;
		16'b0110011011001011: color_data = 12'b001110100111;
		16'b0110011011001100: color_data = 12'b001110100111;
		16'b0110011011001101: color_data = 12'b001110100111;
		16'b0110011011001110: color_data = 12'b001110100111;
		16'b0110011011001111: color_data = 12'b001110100111;
		16'b0110011011010000: color_data = 12'b001110100111;
		16'b0110011011010001: color_data = 12'b001110100111;
		16'b0110011011010010: color_data = 12'b001110100111;
		16'b0110011011010011: color_data = 12'b001110100111;
		16'b0110011011010100: color_data = 12'b001110100111;
		16'b0110011011010101: color_data = 12'b001110100111;
		16'b0110011011010110: color_data = 12'b001110100111;
		16'b0110011011010111: color_data = 12'b001110100111;
		16'b0110011011011000: color_data = 12'b001110100111;
		16'b0110011011011001: color_data = 12'b001110100111;
		16'b0110011011011010: color_data = 12'b001110100111;
		16'b0110011011011011: color_data = 12'b001110100111;
		16'b0110011011011100: color_data = 12'b001110100111;
		16'b0110011011011101: color_data = 12'b001110100111;
		16'b0110011011011110: color_data = 12'b001110100111;
		16'b0110011011011111: color_data = 12'b001110100111;
		16'b0110011011100000: color_data = 12'b001110100111;
		16'b0110011011100001: color_data = 12'b001110100111;
		16'b0110011011100010: color_data = 12'b001110100111;
		16'b0110011011110110: color_data = 12'b001110100111;
		16'b0110011011110111: color_data = 12'b001110100111;
		16'b0110011011111000: color_data = 12'b001110100111;
		16'b0110011011111001: color_data = 12'b001110100111;
		16'b0110011011111010: color_data = 12'b001110100111;
		16'b0110011011111011: color_data = 12'b001110100111;
		16'b0110011011111100: color_data = 12'b001110100111;
		16'b0110011011111101: color_data = 12'b001110100111;
		16'b0110011011111110: color_data = 12'b001110100111;
		16'b0110011011111111: color_data = 12'b001110100111;
		16'b0110011100000000: color_data = 12'b001110100111;
		16'b0110011100000001: color_data = 12'b001110100111;
		16'b0110011100011010: color_data = 12'b001110100111;
		16'b0110011100011011: color_data = 12'b001110100111;
		16'b0110011100011100: color_data = 12'b001110100111;
		16'b0110011100011101: color_data = 12'b001110100111;
		16'b0110011100011110: color_data = 12'b001110100111;
		16'b0110011100011111: color_data = 12'b001110100111;
		16'b0110011100100000: color_data = 12'b001110100111;
		16'b0110011100100001: color_data = 12'b001110100111;
		16'b0110011100100010: color_data = 12'b001110100111;
		16'b0110011100100011: color_data = 12'b001110100111;
		16'b0110011100100100: color_data = 12'b001110100111;
		16'b0110011100100101: color_data = 12'b001110100111;
		16'b0110011100100110: color_data = 12'b001110100111;
		16'b0110011100101101: color_data = 12'b001110100111;
		16'b0110011100101110: color_data = 12'b001110100111;
		16'b0110011100101111: color_data = 12'b001110100111;
		16'b0110011100110000: color_data = 12'b001110100111;
		16'b0110011100110001: color_data = 12'b001110100111;
		16'b0110011100110010: color_data = 12'b001110100111;
		16'b0110011100110011: color_data = 12'b001110100111;
		16'b0110011100110100: color_data = 12'b001110100111;
		16'b0110011100110101: color_data = 12'b001110100111;
		16'b0110011100110110: color_data = 12'b001110100111;
		16'b0110011100110111: color_data = 12'b001110100111;
		16'b0110011100111000: color_data = 12'b001110100111;
		16'b0110011101000101: color_data = 12'b001110100111;
		16'b0110011101000110: color_data = 12'b001110100111;
		16'b0110011101000111: color_data = 12'b001110100111;
		16'b0110011101001000: color_data = 12'b001110100111;
		16'b0110011101001001: color_data = 12'b001110100111;
		16'b0110011101001010: color_data = 12'b001110100111;
		16'b0110011101001011: color_data = 12'b001110100111;
		16'b0110011101001100: color_data = 12'b001110100111;
		16'b0110011101001101: color_data = 12'b001110100111;
		16'b0110011101001110: color_data = 12'b001110100111;
		16'b0110011101001111: color_data = 12'b001110100111;
		16'b0110011101010000: color_data = 12'b001110100111;
		16'b0110011101010001: color_data = 12'b001110100111;
		16'b0110011101011000: color_data = 12'b001110100111;
		16'b0110011101011001: color_data = 12'b001110100111;
		16'b0110011101011010: color_data = 12'b001110100111;
		16'b0110011101011011: color_data = 12'b001110100111;
		16'b0110011101011100: color_data = 12'b001110100111;
		16'b0110011101011101: color_data = 12'b001110100111;
		16'b0110011101011110: color_data = 12'b001110100111;
		16'b0110011101011111: color_data = 12'b001110100111;
		16'b0110011101100000: color_data = 12'b001110100111;
		16'b0110011101100001: color_data = 12'b001110100111;
		16'b0110011101100010: color_data = 12'b001110100111;
		16'b0110011101100011: color_data = 12'b001110100111;
		16'b0110011101110000: color_data = 12'b001110100111;
		16'b0110011101110001: color_data = 12'b001110100111;
		16'b0110011101110010: color_data = 12'b001110100111;
		16'b0110011101110011: color_data = 12'b001110100111;
		16'b0110011101110100: color_data = 12'b001110100111;
		16'b0110011101110101: color_data = 12'b001110100111;
		16'b0110011101110110: color_data = 12'b001110100111;
		16'b0110011101110111: color_data = 12'b001110100111;
		16'b0110011101111000: color_data = 12'b001110100111;
		16'b0110011101111001: color_data = 12'b001110100111;
		16'b0110011101111010: color_data = 12'b001110100111;
		16'b0110011101111011: color_data = 12'b001110100111;
		16'b0110100000000000: color_data = 12'b001110100111;
		16'b0110100000000001: color_data = 12'b001110100111;
		16'b0110100000000010: color_data = 12'b001110100111;
		16'b0110100000000011: color_data = 12'b001110100111;
		16'b0110100000000100: color_data = 12'b001110100111;
		16'b0110100000000101: color_data = 12'b001110100111;
		16'b0110100000000110: color_data = 12'b001110100111;
		16'b0110100000000111: color_data = 12'b001110100111;
		16'b0110100000001000: color_data = 12'b001110100111;
		16'b0110100000001001: color_data = 12'b001110100111;
		16'b0110100000001010: color_data = 12'b001110100111;
		16'b0110100000001011: color_data = 12'b001110100111;
		16'b0110100000001100: color_data = 12'b001110100111;
		16'b0110100000101011: color_data = 12'b001110100111;
		16'b0110100000101100: color_data = 12'b001110100111;
		16'b0110100000101101: color_data = 12'b001110100111;
		16'b0110100000101110: color_data = 12'b001110100111;
		16'b0110100000101111: color_data = 12'b001110100111;
		16'b0110100000110000: color_data = 12'b001110100111;
		16'b0110100000110001: color_data = 12'b001110100111;
		16'b0110100000110010: color_data = 12'b001110100111;
		16'b0110100000110011: color_data = 12'b001110100111;
		16'b0110100000110100: color_data = 12'b001110100111;
		16'b0110100000110101: color_data = 12'b001110100111;
		16'b0110100000110110: color_data = 12'b001110100111;
		16'b0110100000110111: color_data = 12'b001110100111;
		16'b0110100000111000: color_data = 12'b001110100111;
		16'b0110100000111001: color_data = 12'b001110100111;
		16'b0110100000111010: color_data = 12'b001110100111;
		16'b0110100000111011: color_data = 12'b001110100111;
		16'b0110100000111100: color_data = 12'b001110100111;
		16'b0110100000111101: color_data = 12'b001110100111;
		16'b0110100000111110: color_data = 12'b001110100111;
		16'b0110100000111111: color_data = 12'b001110100111;
		16'b0110100001000000: color_data = 12'b001110100111;
		16'b0110100001000001: color_data = 12'b001110100111;
		16'b0110100001000010: color_data = 12'b001110100111;
		16'b0110100001000011: color_data = 12'b001110100111;
		16'b0110100001000100: color_data = 12'b001110100111;
		16'b0110100001000101: color_data = 12'b001110100111;
		16'b0110100001000110: color_data = 12'b001110100111;
		16'b0110100001000111: color_data = 12'b001110100111;
		16'b0110100001001000: color_data = 12'b001110100111;
		16'b0110100001001001: color_data = 12'b001110100111;
		16'b0110100001001010: color_data = 12'b001110100111;
		16'b0110100001001011: color_data = 12'b001110100111;
		16'b0110100001001100: color_data = 12'b001110100111;
		16'b0110100001001101: color_data = 12'b001110100111;
		16'b0110100001001110: color_data = 12'b001110100111;
		16'b0110100001001111: color_data = 12'b001110100111;
		16'b0110100001011100: color_data = 12'b001110100111;
		16'b0110100001011101: color_data = 12'b001110100111;
		16'b0110100001011110: color_data = 12'b001110100111;
		16'b0110100001011111: color_data = 12'b001110100111;
		16'b0110100001100000: color_data = 12'b001110100111;
		16'b0110100001100001: color_data = 12'b001110100111;
		16'b0110100001100010: color_data = 12'b001110100111;
		16'b0110100001100011: color_data = 12'b001110100111;
		16'b0110100001100100: color_data = 12'b001110100111;
		16'b0110100001100101: color_data = 12'b001110100111;
		16'b0110100001100110: color_data = 12'b001110100111;
		16'b0110100001100111: color_data = 12'b001110100111;
		16'b0110100001101000: color_data = 12'b001110100111;
		16'b0110100001110101: color_data = 12'b001110100111;
		16'b0110100001110110: color_data = 12'b001110100111;
		16'b0110100001110111: color_data = 12'b001110100111;
		16'b0110100001111000: color_data = 12'b001110100111;
		16'b0110100001111001: color_data = 12'b001110100111;
		16'b0110100001111010: color_data = 12'b001110100111;
		16'b0110100001111011: color_data = 12'b001110100111;
		16'b0110100001111100: color_data = 12'b001110100111;
		16'b0110100001111101: color_data = 12'b001110100111;
		16'b0110100001111110: color_data = 12'b001110100111;
		16'b0110100001111111: color_data = 12'b001110100111;
		16'b0110100010000000: color_data = 12'b001110100111;
		16'b0110100010001101: color_data = 12'b001110100111;
		16'b0110100010001110: color_data = 12'b001110100111;
		16'b0110100010001111: color_data = 12'b001110100111;
		16'b0110100010010000: color_data = 12'b001110100111;
		16'b0110100010010001: color_data = 12'b001110100111;
		16'b0110100010010010: color_data = 12'b001110100111;
		16'b0110100010010011: color_data = 12'b001110100111;
		16'b0110100010010100: color_data = 12'b001110100111;
		16'b0110100010010101: color_data = 12'b001110100111;
		16'b0110100010010110: color_data = 12'b001110100111;
		16'b0110100010010111: color_data = 12'b001110100111;
		16'b0110100010011000: color_data = 12'b001110100111;
		16'b0110100010011001: color_data = 12'b001110100111;
		16'b0110100010100000: color_data = 12'b001110100111;
		16'b0110100010100001: color_data = 12'b001110100111;
		16'b0110100010100010: color_data = 12'b001110100111;
		16'b0110100010100011: color_data = 12'b001110100111;
		16'b0110100010100100: color_data = 12'b001110100111;
		16'b0110100010100101: color_data = 12'b001110100111;
		16'b0110100010100110: color_data = 12'b001110100111;
		16'b0110100010100111: color_data = 12'b001110100111;
		16'b0110100010101000: color_data = 12'b001110100111;
		16'b0110100010101001: color_data = 12'b001110100111;
		16'b0110100010101010: color_data = 12'b001110100111;
		16'b0110100010101011: color_data = 12'b001110100111;
		16'b0110100010111000: color_data = 12'b001110100111;
		16'b0110100010111001: color_data = 12'b001110100111;
		16'b0110100010111010: color_data = 12'b001110100111;
		16'b0110100010111011: color_data = 12'b001110100111;
		16'b0110100010111100: color_data = 12'b001110100111;
		16'b0110100010111101: color_data = 12'b001110100111;
		16'b0110100010111110: color_data = 12'b001110100111;
		16'b0110100010111111: color_data = 12'b001110100111;
		16'b0110100011000000: color_data = 12'b001110100111;
		16'b0110100011000001: color_data = 12'b001110100111;
		16'b0110100011000010: color_data = 12'b001110100111;
		16'b0110100011000011: color_data = 12'b001110100111;
		16'b0110100011000100: color_data = 12'b001110100111;
		16'b0110100011001011: color_data = 12'b001110100111;
		16'b0110100011001100: color_data = 12'b001110100111;
		16'b0110100011001101: color_data = 12'b001110100111;
		16'b0110100011001110: color_data = 12'b001110100111;
		16'b0110100011001111: color_data = 12'b001110100111;
		16'b0110100011010000: color_data = 12'b001110100111;
		16'b0110100011010001: color_data = 12'b001110100111;
		16'b0110100011010010: color_data = 12'b001110100111;
		16'b0110100011010011: color_data = 12'b001110100111;
		16'b0110100011010100: color_data = 12'b001110100111;
		16'b0110100011010101: color_data = 12'b001110100111;
		16'b0110100011010110: color_data = 12'b001110100111;
		16'b0110100011010111: color_data = 12'b001110100111;
		16'b0110100011011000: color_data = 12'b001110100111;
		16'b0110100011011001: color_data = 12'b001110100111;
		16'b0110100011011010: color_data = 12'b001110100111;
		16'b0110100011011011: color_data = 12'b001110100111;
		16'b0110100011011100: color_data = 12'b001110100111;
		16'b0110100011011101: color_data = 12'b001110100111;
		16'b0110100011011110: color_data = 12'b001110100111;
		16'b0110100011011111: color_data = 12'b001110100111;
		16'b0110100011100000: color_data = 12'b001110100111;
		16'b0110100011100001: color_data = 12'b001110100111;
		16'b0110100011100010: color_data = 12'b001110100111;
		16'b0110100011110110: color_data = 12'b001110100111;
		16'b0110100011110111: color_data = 12'b001110100111;
		16'b0110100011111000: color_data = 12'b001110100111;
		16'b0110100011111001: color_data = 12'b001110100111;
		16'b0110100011111010: color_data = 12'b001110100111;
		16'b0110100011111011: color_data = 12'b001110100111;
		16'b0110100011111100: color_data = 12'b001110100111;
		16'b0110100011111101: color_data = 12'b001110100111;
		16'b0110100011111110: color_data = 12'b001110100111;
		16'b0110100011111111: color_data = 12'b001110100111;
		16'b0110100100000000: color_data = 12'b001110100111;
		16'b0110100100000001: color_data = 12'b001110100111;
		16'b0110100100011010: color_data = 12'b001110100111;
		16'b0110100100011011: color_data = 12'b001110100111;
		16'b0110100100011100: color_data = 12'b001110100111;
		16'b0110100100011101: color_data = 12'b001110100111;
		16'b0110100100011110: color_data = 12'b001110100111;
		16'b0110100100011111: color_data = 12'b001110100111;
		16'b0110100100100000: color_data = 12'b001110100111;
		16'b0110100100100001: color_data = 12'b001110100111;
		16'b0110100100100010: color_data = 12'b001110100111;
		16'b0110100100100011: color_data = 12'b001110100111;
		16'b0110100100100100: color_data = 12'b001110100111;
		16'b0110100100100101: color_data = 12'b001110100111;
		16'b0110100100100110: color_data = 12'b001110100111;
		16'b0110100100101101: color_data = 12'b001110100111;
		16'b0110100100101110: color_data = 12'b001110100111;
		16'b0110100100101111: color_data = 12'b001110100111;
		16'b0110100100110000: color_data = 12'b001110100111;
		16'b0110100100110001: color_data = 12'b001110100111;
		16'b0110100100110010: color_data = 12'b001110100111;
		16'b0110100100110011: color_data = 12'b001110100111;
		16'b0110100100110100: color_data = 12'b001110100111;
		16'b0110100100110101: color_data = 12'b001110100111;
		16'b0110100100110110: color_data = 12'b001110100111;
		16'b0110100100110111: color_data = 12'b001110100111;
		16'b0110100100111000: color_data = 12'b001110100111;
		16'b0110100101000101: color_data = 12'b001110100111;
		16'b0110100101000110: color_data = 12'b001110100111;
		16'b0110100101000111: color_data = 12'b001110100111;
		16'b0110100101001000: color_data = 12'b001110100111;
		16'b0110100101001001: color_data = 12'b001110100111;
		16'b0110100101001010: color_data = 12'b001110100111;
		16'b0110100101001011: color_data = 12'b001110100111;
		16'b0110100101001100: color_data = 12'b001110100111;
		16'b0110100101001101: color_data = 12'b001110100111;
		16'b0110100101001110: color_data = 12'b001110100111;
		16'b0110100101001111: color_data = 12'b001110100111;
		16'b0110100101010000: color_data = 12'b001110100111;
		16'b0110100101010001: color_data = 12'b001110100111;
		16'b0110100101011000: color_data = 12'b001110100111;
		16'b0110100101011001: color_data = 12'b001110100111;
		16'b0110100101011010: color_data = 12'b001110100111;
		16'b0110100101011011: color_data = 12'b001110100111;
		16'b0110100101011100: color_data = 12'b001110100111;
		16'b0110100101011101: color_data = 12'b001110100111;
		16'b0110100101011110: color_data = 12'b001110100111;
		16'b0110100101011111: color_data = 12'b001110100111;
		16'b0110100101100000: color_data = 12'b001110100111;
		16'b0110100101100001: color_data = 12'b001110100111;
		16'b0110100101100010: color_data = 12'b001110100111;
		16'b0110100101100011: color_data = 12'b001110100111;
		16'b0110100101110000: color_data = 12'b001110100111;
		16'b0110100101110001: color_data = 12'b001110100111;
		16'b0110100101110010: color_data = 12'b001110100111;
		16'b0110100101110011: color_data = 12'b001110100111;
		16'b0110100101110100: color_data = 12'b001110100111;
		16'b0110100101110101: color_data = 12'b001110100111;
		16'b0110100101110110: color_data = 12'b001110100111;
		16'b0110100101110111: color_data = 12'b001110100111;
		16'b0110100101111000: color_data = 12'b001110100111;
		16'b0110100101111001: color_data = 12'b001110100111;
		16'b0110100101111010: color_data = 12'b001110100111;
		16'b0110100101111011: color_data = 12'b001110100111;
		16'b0110101000000000: color_data = 12'b001110100111;
		16'b0110101000000001: color_data = 12'b001110100111;
		16'b0110101000000010: color_data = 12'b001110100111;
		16'b0110101000000011: color_data = 12'b001110100111;
		16'b0110101000000100: color_data = 12'b001110100111;
		16'b0110101000000101: color_data = 12'b001110100111;
		16'b0110101000000110: color_data = 12'b001110100111;
		16'b0110101000000111: color_data = 12'b001110100111;
		16'b0110101000001000: color_data = 12'b001110100111;
		16'b0110101000001001: color_data = 12'b001110100111;
		16'b0110101000001010: color_data = 12'b001110100111;
		16'b0110101000001011: color_data = 12'b001110100111;
		16'b0110101000001100: color_data = 12'b001110100111;
		16'b0110101000101011: color_data = 12'b001110100111;
		16'b0110101000101100: color_data = 12'b001110100111;
		16'b0110101000101101: color_data = 12'b001110100111;
		16'b0110101000101110: color_data = 12'b001110100111;
		16'b0110101000101111: color_data = 12'b001110100111;
		16'b0110101000110000: color_data = 12'b001110100111;
		16'b0110101000110001: color_data = 12'b001110100111;
		16'b0110101000110010: color_data = 12'b001110100111;
		16'b0110101000110011: color_data = 12'b001110100111;
		16'b0110101000110100: color_data = 12'b001110100111;
		16'b0110101000110101: color_data = 12'b001110100111;
		16'b0110101000110110: color_data = 12'b001110100111;
		16'b0110101000110111: color_data = 12'b001110100111;
		16'b0110101000111000: color_data = 12'b001110100111;
		16'b0110101000111001: color_data = 12'b001110100111;
		16'b0110101000111010: color_data = 12'b001110100111;
		16'b0110101000111011: color_data = 12'b001110100111;
		16'b0110101000111100: color_data = 12'b001110100111;
		16'b0110101000111101: color_data = 12'b001110100111;
		16'b0110101000111110: color_data = 12'b001110100111;
		16'b0110101000111111: color_data = 12'b001110100111;
		16'b0110101001000000: color_data = 12'b001110100111;
		16'b0110101001000001: color_data = 12'b001110100111;
		16'b0110101001000010: color_data = 12'b001110100111;
		16'b0110101001000011: color_data = 12'b001110100111;
		16'b0110101001000100: color_data = 12'b001110100111;
		16'b0110101001000101: color_data = 12'b001110100111;
		16'b0110101001000110: color_data = 12'b001110100111;
		16'b0110101001000111: color_data = 12'b001110100111;
		16'b0110101001001000: color_data = 12'b001110100111;
		16'b0110101001001001: color_data = 12'b001110100111;
		16'b0110101001001010: color_data = 12'b001110100111;
		16'b0110101001001011: color_data = 12'b001110100111;
		16'b0110101001001100: color_data = 12'b001110100111;
		16'b0110101001001101: color_data = 12'b001110100111;
		16'b0110101001001110: color_data = 12'b001110100111;
		16'b0110101001001111: color_data = 12'b001110100111;
		16'b0110101001011100: color_data = 12'b001110100111;
		16'b0110101001011101: color_data = 12'b001110100111;
		16'b0110101001011110: color_data = 12'b001110100111;
		16'b0110101001011111: color_data = 12'b001110100111;
		16'b0110101001100000: color_data = 12'b001110100111;
		16'b0110101001100001: color_data = 12'b001110100111;
		16'b0110101001100010: color_data = 12'b001110100111;
		16'b0110101001100011: color_data = 12'b001110100111;
		16'b0110101001100100: color_data = 12'b001110100111;
		16'b0110101001100101: color_data = 12'b001110100111;
		16'b0110101001100110: color_data = 12'b001110100111;
		16'b0110101001100111: color_data = 12'b001110100111;
		16'b0110101001101000: color_data = 12'b001110100111;
		16'b0110101001110101: color_data = 12'b001110100111;
		16'b0110101001110110: color_data = 12'b001110100111;
		16'b0110101001110111: color_data = 12'b001110100111;
		16'b0110101001111000: color_data = 12'b001110100111;
		16'b0110101001111001: color_data = 12'b001110100111;
		16'b0110101001111010: color_data = 12'b001110100111;
		16'b0110101001111011: color_data = 12'b001110100111;
		16'b0110101001111100: color_data = 12'b001110100111;
		16'b0110101001111101: color_data = 12'b001110100111;
		16'b0110101001111110: color_data = 12'b001110100111;
		16'b0110101001111111: color_data = 12'b001110100111;
		16'b0110101010000000: color_data = 12'b001110100111;
		16'b0110101010001101: color_data = 12'b001110100111;
		16'b0110101010001110: color_data = 12'b001110100111;
		16'b0110101010001111: color_data = 12'b001110100111;
		16'b0110101010010000: color_data = 12'b001110100111;
		16'b0110101010010001: color_data = 12'b001110100111;
		16'b0110101010010010: color_data = 12'b001110100111;
		16'b0110101010010011: color_data = 12'b001110100111;
		16'b0110101010010100: color_data = 12'b001110100111;
		16'b0110101010010101: color_data = 12'b001110100111;
		16'b0110101010010110: color_data = 12'b001110100111;
		16'b0110101010010111: color_data = 12'b001110100111;
		16'b0110101010011000: color_data = 12'b001110100111;
		16'b0110101010011001: color_data = 12'b001110100111;
		16'b0110101010100000: color_data = 12'b001110100111;
		16'b0110101010100001: color_data = 12'b001110100111;
		16'b0110101010100010: color_data = 12'b001110100111;
		16'b0110101010100011: color_data = 12'b001110100111;
		16'b0110101010100100: color_data = 12'b001110100111;
		16'b0110101010100101: color_data = 12'b001110100111;
		16'b0110101010100110: color_data = 12'b001110100111;
		16'b0110101010100111: color_data = 12'b001110100111;
		16'b0110101010101000: color_data = 12'b001110100111;
		16'b0110101010101001: color_data = 12'b001110100111;
		16'b0110101010101010: color_data = 12'b001110100111;
		16'b0110101010101011: color_data = 12'b001110100111;
		16'b0110101010111000: color_data = 12'b001110100111;
		16'b0110101010111001: color_data = 12'b001110100111;
		16'b0110101010111010: color_data = 12'b001110100111;
		16'b0110101010111011: color_data = 12'b001110100111;
		16'b0110101010111100: color_data = 12'b001110100111;
		16'b0110101010111101: color_data = 12'b001110100111;
		16'b0110101010111110: color_data = 12'b001110100111;
		16'b0110101010111111: color_data = 12'b001110100111;
		16'b0110101011000000: color_data = 12'b001110100111;
		16'b0110101011000001: color_data = 12'b001110100111;
		16'b0110101011000010: color_data = 12'b001110100111;
		16'b0110101011000011: color_data = 12'b001110100111;
		16'b0110101011000100: color_data = 12'b001110100111;
		16'b0110101011001011: color_data = 12'b001110100111;
		16'b0110101011001100: color_data = 12'b001110100111;
		16'b0110101011001101: color_data = 12'b001110100111;
		16'b0110101011001110: color_data = 12'b001110100111;
		16'b0110101011001111: color_data = 12'b001110100111;
		16'b0110101011010000: color_data = 12'b001110100111;
		16'b0110101011010001: color_data = 12'b001110100111;
		16'b0110101011010010: color_data = 12'b001110100111;
		16'b0110101011010011: color_data = 12'b001110100111;
		16'b0110101011010100: color_data = 12'b001110100111;
		16'b0110101011010101: color_data = 12'b001110100111;
		16'b0110101011010110: color_data = 12'b001110100111;
		16'b0110101011010111: color_data = 12'b001110100111;
		16'b0110101011011000: color_data = 12'b001110100111;
		16'b0110101011011001: color_data = 12'b001110100111;
		16'b0110101011011010: color_data = 12'b001110100111;
		16'b0110101011011011: color_data = 12'b001110100111;
		16'b0110101011011100: color_data = 12'b001110100111;
		16'b0110101011011101: color_data = 12'b001110100111;
		16'b0110101011011110: color_data = 12'b001110100111;
		16'b0110101011011111: color_data = 12'b001110100111;
		16'b0110101011100000: color_data = 12'b001110100111;
		16'b0110101011100001: color_data = 12'b001110100111;
		16'b0110101011100010: color_data = 12'b001110100111;
		16'b0110101011110110: color_data = 12'b001110100111;
		16'b0110101011110111: color_data = 12'b001110100111;
		16'b0110101011111000: color_data = 12'b001110100111;
		16'b0110101011111001: color_data = 12'b001110100111;
		16'b0110101011111010: color_data = 12'b001110100111;
		16'b0110101011111011: color_data = 12'b001110100111;
		16'b0110101011111100: color_data = 12'b001110100111;
		16'b0110101011111101: color_data = 12'b001110100111;
		16'b0110101011111110: color_data = 12'b001110100111;
		16'b0110101011111111: color_data = 12'b001110100111;
		16'b0110101100000000: color_data = 12'b001110100111;
		16'b0110101100000001: color_data = 12'b001110100111;
		16'b0110101100011010: color_data = 12'b001110100111;
		16'b0110101100011011: color_data = 12'b001110100111;
		16'b0110101100011100: color_data = 12'b001110100111;
		16'b0110101100011101: color_data = 12'b001110100111;
		16'b0110101100011110: color_data = 12'b001110100111;
		16'b0110101100011111: color_data = 12'b001110100111;
		16'b0110101100100000: color_data = 12'b001110100111;
		16'b0110101100100001: color_data = 12'b001110100111;
		16'b0110101100100010: color_data = 12'b001110100111;
		16'b0110101100100011: color_data = 12'b001110100111;
		16'b0110101100100100: color_data = 12'b001110100111;
		16'b0110101100100101: color_data = 12'b001110100111;
		16'b0110101100100110: color_data = 12'b001110100111;
		16'b0110101100101101: color_data = 12'b001110100111;
		16'b0110101100101110: color_data = 12'b001110100111;
		16'b0110101100101111: color_data = 12'b001110100111;
		16'b0110101100110000: color_data = 12'b001110100111;
		16'b0110101100110001: color_data = 12'b001110100111;
		16'b0110101100110010: color_data = 12'b001110100111;
		16'b0110101100110011: color_data = 12'b001110100111;
		16'b0110101100110100: color_data = 12'b001110100111;
		16'b0110101100110101: color_data = 12'b001110100111;
		16'b0110101100110110: color_data = 12'b001110100111;
		16'b0110101100110111: color_data = 12'b001110100111;
		16'b0110101100111000: color_data = 12'b001110100111;
		16'b0110101101000101: color_data = 12'b001110100111;
		16'b0110101101000110: color_data = 12'b001110100111;
		16'b0110101101000111: color_data = 12'b001110100111;
		16'b0110101101001000: color_data = 12'b001110100111;
		16'b0110101101001001: color_data = 12'b001110100111;
		16'b0110101101001010: color_data = 12'b001110100111;
		16'b0110101101001011: color_data = 12'b001110100111;
		16'b0110101101001100: color_data = 12'b001110100111;
		16'b0110101101001101: color_data = 12'b001110100111;
		16'b0110101101001110: color_data = 12'b001110100111;
		16'b0110101101001111: color_data = 12'b001110100111;
		16'b0110101101010000: color_data = 12'b001110100111;
		16'b0110101101010001: color_data = 12'b001110100111;
		16'b0110101101011000: color_data = 12'b001110100111;
		16'b0110101101011001: color_data = 12'b001110100111;
		16'b0110101101011010: color_data = 12'b001110100111;
		16'b0110101101011011: color_data = 12'b001110100111;
		16'b0110101101011100: color_data = 12'b001110100111;
		16'b0110101101011101: color_data = 12'b001110100111;
		16'b0110101101011110: color_data = 12'b001110100111;
		16'b0110101101011111: color_data = 12'b001110100111;
		16'b0110101101100000: color_data = 12'b001110100111;
		16'b0110101101100001: color_data = 12'b001110100111;
		16'b0110101101100010: color_data = 12'b001110100111;
		16'b0110101101100011: color_data = 12'b001110100111;
		16'b0110101101110000: color_data = 12'b001110100111;
		16'b0110101101110001: color_data = 12'b001110100111;
		16'b0110101101110010: color_data = 12'b001110100111;
		16'b0110101101110011: color_data = 12'b001110100111;
		16'b0110101101110100: color_data = 12'b001110100111;
		16'b0110101101110101: color_data = 12'b001110100111;
		16'b0110101101110110: color_data = 12'b001110100111;
		16'b0110101101110111: color_data = 12'b001110100111;
		16'b0110101101111000: color_data = 12'b001110100111;
		16'b0110101101111001: color_data = 12'b001110100111;
		16'b0110101101111010: color_data = 12'b001110100111;
		16'b0110101101111011: color_data = 12'b001110100111;
		16'b0110110000000000: color_data = 12'b001110100111;
		16'b0110110000000001: color_data = 12'b001110100111;
		16'b0110110000000010: color_data = 12'b001110100111;
		16'b0110110000000011: color_data = 12'b001110100111;
		16'b0110110000000100: color_data = 12'b001110100111;
		16'b0110110000000101: color_data = 12'b001110100111;
		16'b0110110000000110: color_data = 12'b001110100111;
		16'b0110110000000111: color_data = 12'b001110100111;
		16'b0110110000001000: color_data = 12'b001110100111;
		16'b0110110000001001: color_data = 12'b001110100111;
		16'b0110110000001010: color_data = 12'b001110100111;
		16'b0110110000001011: color_data = 12'b001110100111;
		16'b0110110000001100: color_data = 12'b001110100111;
		16'b0110110000101011: color_data = 12'b001110100111;
		16'b0110110000101100: color_data = 12'b001110100111;
		16'b0110110000101101: color_data = 12'b001110100111;
		16'b0110110000101110: color_data = 12'b001110100111;
		16'b0110110000101111: color_data = 12'b001110100111;
		16'b0110110000110000: color_data = 12'b001110100111;
		16'b0110110000110001: color_data = 12'b001110100111;
		16'b0110110000110010: color_data = 12'b001110100111;
		16'b0110110000110011: color_data = 12'b001110100111;
		16'b0110110000110100: color_data = 12'b001110100111;
		16'b0110110000110101: color_data = 12'b001110100111;
		16'b0110110000110110: color_data = 12'b001110100111;
		16'b0110110000110111: color_data = 12'b001110100111;
		16'b0110110000111000: color_data = 12'b001110100111;
		16'b0110110000111001: color_data = 12'b001110100111;
		16'b0110110000111010: color_data = 12'b001110100111;
		16'b0110110000111011: color_data = 12'b001110100111;
		16'b0110110000111100: color_data = 12'b001110100111;
		16'b0110110000111101: color_data = 12'b001110100111;
		16'b0110110000111110: color_data = 12'b001110100111;
		16'b0110110000111111: color_data = 12'b001110100111;
		16'b0110110001000000: color_data = 12'b001110100111;
		16'b0110110001000001: color_data = 12'b001110100111;
		16'b0110110001000010: color_data = 12'b001110100111;
		16'b0110110001000011: color_data = 12'b001110100111;
		16'b0110110001000100: color_data = 12'b001110100111;
		16'b0110110001000101: color_data = 12'b001110100111;
		16'b0110110001000110: color_data = 12'b001110100111;
		16'b0110110001000111: color_data = 12'b001110100111;
		16'b0110110001001000: color_data = 12'b001110100111;
		16'b0110110001001001: color_data = 12'b001110100111;
		16'b0110110001001010: color_data = 12'b001110100111;
		16'b0110110001001011: color_data = 12'b001110100111;
		16'b0110110001001100: color_data = 12'b001110100111;
		16'b0110110001001101: color_data = 12'b001110100111;
		16'b0110110001001110: color_data = 12'b001110100111;
		16'b0110110001001111: color_data = 12'b001110100111;
		16'b0110110001011100: color_data = 12'b001110100111;
		16'b0110110001011101: color_data = 12'b001110100111;
		16'b0110110001011110: color_data = 12'b001110100111;
		16'b0110110001011111: color_data = 12'b001110100111;
		16'b0110110001100000: color_data = 12'b001110100111;
		16'b0110110001100001: color_data = 12'b001110100111;
		16'b0110110001100010: color_data = 12'b001110100111;
		16'b0110110001100011: color_data = 12'b001110100111;
		16'b0110110001100100: color_data = 12'b001110100111;
		16'b0110110001100101: color_data = 12'b001110100111;
		16'b0110110001100110: color_data = 12'b001110100111;
		16'b0110110001100111: color_data = 12'b001110100111;
		16'b0110110001101000: color_data = 12'b001110100111;
		16'b0110110001110101: color_data = 12'b001110100111;
		16'b0110110001110110: color_data = 12'b001110100111;
		16'b0110110001110111: color_data = 12'b001110100111;
		16'b0110110001111000: color_data = 12'b001110100111;
		16'b0110110001111001: color_data = 12'b001110100111;
		16'b0110110001111010: color_data = 12'b001110100111;
		16'b0110110001111011: color_data = 12'b001110100111;
		16'b0110110001111100: color_data = 12'b001110100111;
		16'b0110110001111101: color_data = 12'b001110100111;
		16'b0110110001111110: color_data = 12'b001110100111;
		16'b0110110001111111: color_data = 12'b001110100111;
		16'b0110110010000000: color_data = 12'b001110100111;
		16'b0110110010001101: color_data = 12'b001110100111;
		16'b0110110010001110: color_data = 12'b001110100111;
		16'b0110110010001111: color_data = 12'b001110100111;
		16'b0110110010010000: color_data = 12'b001110100111;
		16'b0110110010010001: color_data = 12'b001110100111;
		16'b0110110010010010: color_data = 12'b001110100111;
		16'b0110110010010011: color_data = 12'b001110100111;
		16'b0110110010010100: color_data = 12'b001110100111;
		16'b0110110010010101: color_data = 12'b001110100111;
		16'b0110110010010110: color_data = 12'b001110100111;
		16'b0110110010010111: color_data = 12'b001110100111;
		16'b0110110010011000: color_data = 12'b001110100111;
		16'b0110110010011001: color_data = 12'b001110100111;
		16'b0110110010100000: color_data = 12'b001110100111;
		16'b0110110010100001: color_data = 12'b001110100111;
		16'b0110110010100010: color_data = 12'b001110100111;
		16'b0110110010100011: color_data = 12'b001110100111;
		16'b0110110010100100: color_data = 12'b001110100111;
		16'b0110110010100101: color_data = 12'b001110100111;
		16'b0110110010100110: color_data = 12'b001110100111;
		16'b0110110010100111: color_data = 12'b001110100111;
		16'b0110110010101000: color_data = 12'b001110100111;
		16'b0110110010101001: color_data = 12'b001110100111;
		16'b0110110010101010: color_data = 12'b001110100111;
		16'b0110110010101011: color_data = 12'b001110100111;
		16'b0110110010111000: color_data = 12'b001110100111;
		16'b0110110010111001: color_data = 12'b001110100111;
		16'b0110110010111010: color_data = 12'b001110100111;
		16'b0110110010111011: color_data = 12'b001110100111;
		16'b0110110010111100: color_data = 12'b001110100111;
		16'b0110110010111101: color_data = 12'b001110100111;
		16'b0110110010111110: color_data = 12'b001110100111;
		16'b0110110010111111: color_data = 12'b001110100111;
		16'b0110110011000000: color_data = 12'b001110100111;
		16'b0110110011000001: color_data = 12'b001110100111;
		16'b0110110011000010: color_data = 12'b001110100111;
		16'b0110110011000011: color_data = 12'b001110100111;
		16'b0110110011000100: color_data = 12'b001110100111;
		16'b0110110011001011: color_data = 12'b001110100111;
		16'b0110110011001100: color_data = 12'b001110100111;
		16'b0110110011001101: color_data = 12'b001110100111;
		16'b0110110011001110: color_data = 12'b001110100111;
		16'b0110110011001111: color_data = 12'b001110100111;
		16'b0110110011010000: color_data = 12'b001110100111;
		16'b0110110011010001: color_data = 12'b001110100111;
		16'b0110110011010010: color_data = 12'b001110100111;
		16'b0110110011010011: color_data = 12'b001110100111;
		16'b0110110011010100: color_data = 12'b001110100111;
		16'b0110110011010101: color_data = 12'b001110100111;
		16'b0110110011010110: color_data = 12'b001110100111;
		16'b0110110011010111: color_data = 12'b001110100111;
		16'b0110110011011000: color_data = 12'b001110100111;
		16'b0110110011011001: color_data = 12'b001110100111;
		16'b0110110011011010: color_data = 12'b001110100111;
		16'b0110110011011011: color_data = 12'b001110100111;
		16'b0110110011011100: color_data = 12'b001110100111;
		16'b0110110011011101: color_data = 12'b001110100111;
		16'b0110110011011110: color_data = 12'b001110100111;
		16'b0110110011011111: color_data = 12'b001110100111;
		16'b0110110011100000: color_data = 12'b001110100111;
		16'b0110110011100001: color_data = 12'b001110100111;
		16'b0110110011100010: color_data = 12'b001110100111;
		16'b0110110011110110: color_data = 12'b001110100111;
		16'b0110110011110111: color_data = 12'b001110100111;
		16'b0110110011111000: color_data = 12'b001110100111;
		16'b0110110011111001: color_data = 12'b001110100111;
		16'b0110110011111010: color_data = 12'b001110100111;
		16'b0110110011111011: color_data = 12'b001110100111;
		16'b0110110011111100: color_data = 12'b001110100111;
		16'b0110110011111101: color_data = 12'b001110100111;
		16'b0110110011111110: color_data = 12'b001110100111;
		16'b0110110011111111: color_data = 12'b001110100111;
		16'b0110110100000000: color_data = 12'b001110100111;
		16'b0110110100000001: color_data = 12'b001110100111;
		16'b0110110100011010: color_data = 12'b001110100111;
		16'b0110110100011011: color_data = 12'b001110100111;
		16'b0110110100011100: color_data = 12'b001110100111;
		16'b0110110100011101: color_data = 12'b001110100111;
		16'b0110110100011110: color_data = 12'b001110100111;
		16'b0110110100011111: color_data = 12'b001110100111;
		16'b0110110100100000: color_data = 12'b001110100111;
		16'b0110110100100001: color_data = 12'b001110100111;
		16'b0110110100100010: color_data = 12'b001110100111;
		16'b0110110100100011: color_data = 12'b001110100111;
		16'b0110110100100100: color_data = 12'b001110100111;
		16'b0110110100100101: color_data = 12'b001110100111;
		16'b0110110100100110: color_data = 12'b001110100111;
		16'b0110110100101101: color_data = 12'b001110100111;
		16'b0110110100101110: color_data = 12'b001110100111;
		16'b0110110100101111: color_data = 12'b001110100111;
		16'b0110110100110000: color_data = 12'b001110100111;
		16'b0110110100110001: color_data = 12'b001110100111;
		16'b0110110100110010: color_data = 12'b001110100111;
		16'b0110110100110011: color_data = 12'b001110100111;
		16'b0110110100110100: color_data = 12'b001110100111;
		16'b0110110100110101: color_data = 12'b001110100111;
		16'b0110110100110110: color_data = 12'b001110100111;
		16'b0110110100110111: color_data = 12'b001110100111;
		16'b0110110100111000: color_data = 12'b001110100111;
		16'b0110110101000101: color_data = 12'b001110100111;
		16'b0110110101000110: color_data = 12'b001110100111;
		16'b0110110101000111: color_data = 12'b001110100111;
		16'b0110110101001000: color_data = 12'b001110100111;
		16'b0110110101001001: color_data = 12'b001110100111;
		16'b0110110101001010: color_data = 12'b001110100111;
		16'b0110110101001011: color_data = 12'b001110100111;
		16'b0110110101001100: color_data = 12'b001110100111;
		16'b0110110101001101: color_data = 12'b001110100111;
		16'b0110110101001110: color_data = 12'b001110100111;
		16'b0110110101001111: color_data = 12'b001110100111;
		16'b0110110101010000: color_data = 12'b001110100111;
		16'b0110110101010001: color_data = 12'b001110100111;
		16'b0110110101011000: color_data = 12'b001110100111;
		16'b0110110101011001: color_data = 12'b001110100111;
		16'b0110110101011010: color_data = 12'b001110100111;
		16'b0110110101011011: color_data = 12'b001110100111;
		16'b0110110101011100: color_data = 12'b001110100111;
		16'b0110110101011101: color_data = 12'b001110100111;
		16'b0110110101011110: color_data = 12'b001110100111;
		16'b0110110101011111: color_data = 12'b001110100111;
		16'b0110110101100000: color_data = 12'b001110100111;
		16'b0110110101100001: color_data = 12'b001110100111;
		16'b0110110101100010: color_data = 12'b001110100111;
		16'b0110110101100011: color_data = 12'b001110100111;
		16'b0110110101110000: color_data = 12'b001110100111;
		16'b0110110101110001: color_data = 12'b001110100111;
		16'b0110110101110010: color_data = 12'b001110100111;
		16'b0110110101110011: color_data = 12'b001110100111;
		16'b0110110101110100: color_data = 12'b001110100111;
		16'b0110110101110101: color_data = 12'b001110100111;
		16'b0110110101110110: color_data = 12'b001110100111;
		16'b0110110101110111: color_data = 12'b001110100111;
		16'b0110110101111000: color_data = 12'b001110100111;
		16'b0110110101111001: color_data = 12'b001110100111;
		16'b0110110101111010: color_data = 12'b001110100111;
		16'b0110110101111011: color_data = 12'b001110100111;
		16'b0110111000000000: color_data = 12'b001110100111;
		16'b0110111000000001: color_data = 12'b001110100111;
		16'b0110111000000010: color_data = 12'b001110100111;
		16'b0110111000000011: color_data = 12'b001110100111;
		16'b0110111000000100: color_data = 12'b001110100111;
		16'b0110111000000101: color_data = 12'b001110100111;
		16'b0110111000000110: color_data = 12'b001110100111;
		16'b0110111000000111: color_data = 12'b001110100111;
		16'b0110111000001000: color_data = 12'b001110100111;
		16'b0110111000001001: color_data = 12'b001110100111;
		16'b0110111000001010: color_data = 12'b001110100111;
		16'b0110111000001011: color_data = 12'b001110100111;
		16'b0110111000001100: color_data = 12'b001110100111;
		16'b0110111000101011: color_data = 12'b001110100111;
		16'b0110111000101100: color_data = 12'b001110100111;
		16'b0110111000101101: color_data = 12'b001110100111;
		16'b0110111000101110: color_data = 12'b001110100111;
		16'b0110111000101111: color_data = 12'b001110100111;
		16'b0110111000110000: color_data = 12'b001110100111;
		16'b0110111000110001: color_data = 12'b001110100111;
		16'b0110111000110010: color_data = 12'b001110100111;
		16'b0110111000110011: color_data = 12'b001110100111;
		16'b0110111000110100: color_data = 12'b001110100111;
		16'b0110111000110101: color_data = 12'b001110100111;
		16'b0110111000110110: color_data = 12'b001110100111;
		16'b0110111000110111: color_data = 12'b001110100111;
		16'b0110111000111000: color_data = 12'b001110100111;
		16'b0110111000111001: color_data = 12'b001110100111;
		16'b0110111000111010: color_data = 12'b001110100111;
		16'b0110111000111011: color_data = 12'b001110100111;
		16'b0110111000111100: color_data = 12'b001110100111;
		16'b0110111000111101: color_data = 12'b001110100111;
		16'b0110111000111110: color_data = 12'b001110100111;
		16'b0110111000111111: color_data = 12'b001110100111;
		16'b0110111001000000: color_data = 12'b001110100111;
		16'b0110111001000001: color_data = 12'b001110100111;
		16'b0110111001000010: color_data = 12'b001110100111;
		16'b0110111001000011: color_data = 12'b001110100111;
		16'b0110111001000100: color_data = 12'b001110100111;
		16'b0110111001000101: color_data = 12'b001110100111;
		16'b0110111001000110: color_data = 12'b001110100111;
		16'b0110111001000111: color_data = 12'b001110100111;
		16'b0110111001001000: color_data = 12'b001110100111;
		16'b0110111001001001: color_data = 12'b001110100111;
		16'b0110111001001010: color_data = 12'b001110100111;
		16'b0110111001001011: color_data = 12'b001110100111;
		16'b0110111001001100: color_data = 12'b001110100111;
		16'b0110111001001101: color_data = 12'b001110100111;
		16'b0110111001001110: color_data = 12'b001110100111;
		16'b0110111001001111: color_data = 12'b001110100111;
		16'b0110111001011100: color_data = 12'b001110100111;
		16'b0110111001011101: color_data = 12'b001110100111;
		16'b0110111001011110: color_data = 12'b001110100111;
		16'b0110111001011111: color_data = 12'b001110100111;
		16'b0110111001100000: color_data = 12'b001110100111;
		16'b0110111001100001: color_data = 12'b001110100111;
		16'b0110111001100010: color_data = 12'b001110100111;
		16'b0110111001100011: color_data = 12'b001110100111;
		16'b0110111001100100: color_data = 12'b001110100111;
		16'b0110111001100101: color_data = 12'b001110100111;
		16'b0110111001100110: color_data = 12'b001110100111;
		16'b0110111001100111: color_data = 12'b001110100111;
		16'b0110111001101000: color_data = 12'b001110100111;
		16'b0110111001110101: color_data = 12'b001110100111;
		16'b0110111001110110: color_data = 12'b001110100111;
		16'b0110111001110111: color_data = 12'b001110100111;
		16'b0110111001111000: color_data = 12'b001110100111;
		16'b0110111001111001: color_data = 12'b001110100111;
		16'b0110111001111010: color_data = 12'b001110100111;
		16'b0110111001111011: color_data = 12'b001110100111;
		16'b0110111001111100: color_data = 12'b001110100111;
		16'b0110111001111101: color_data = 12'b001110100111;
		16'b0110111001111110: color_data = 12'b001110100111;
		16'b0110111001111111: color_data = 12'b001110100111;
		16'b0110111010000000: color_data = 12'b001110100111;
		16'b0110111010001101: color_data = 12'b001110100111;
		16'b0110111010001110: color_data = 12'b001110100111;
		16'b0110111010001111: color_data = 12'b001110100111;
		16'b0110111010010000: color_data = 12'b001110100111;
		16'b0110111010010001: color_data = 12'b001110100111;
		16'b0110111010010010: color_data = 12'b001110100111;
		16'b0110111010010011: color_data = 12'b001110100111;
		16'b0110111010010100: color_data = 12'b001110100111;
		16'b0110111010010101: color_data = 12'b001110100111;
		16'b0110111010010110: color_data = 12'b001110100111;
		16'b0110111010010111: color_data = 12'b001110100111;
		16'b0110111010011000: color_data = 12'b001110100111;
		16'b0110111010011001: color_data = 12'b001110100111;
		16'b0110111010100000: color_data = 12'b001110100111;
		16'b0110111010100001: color_data = 12'b001110100111;
		16'b0110111010100010: color_data = 12'b001110100111;
		16'b0110111010100011: color_data = 12'b001110100111;
		16'b0110111010100100: color_data = 12'b001110100111;
		16'b0110111010100101: color_data = 12'b001110100111;
		16'b0110111010100110: color_data = 12'b001110100111;
		16'b0110111010100111: color_data = 12'b001110100111;
		16'b0110111010101000: color_data = 12'b001110100111;
		16'b0110111010101001: color_data = 12'b001110100111;
		16'b0110111010101010: color_data = 12'b001110100111;
		16'b0110111010101011: color_data = 12'b001110100111;
		16'b0110111010111000: color_data = 12'b001110100111;
		16'b0110111010111001: color_data = 12'b001110100111;
		16'b0110111010111010: color_data = 12'b001110100111;
		16'b0110111010111011: color_data = 12'b001110100111;
		16'b0110111010111100: color_data = 12'b001110100111;
		16'b0110111010111101: color_data = 12'b001110100111;
		16'b0110111010111110: color_data = 12'b001110100111;
		16'b0110111010111111: color_data = 12'b001110100111;
		16'b0110111011000000: color_data = 12'b001110100111;
		16'b0110111011000001: color_data = 12'b001110100111;
		16'b0110111011000010: color_data = 12'b001110100111;
		16'b0110111011000011: color_data = 12'b001110100111;
		16'b0110111011000100: color_data = 12'b001110100111;
		16'b0110111011001011: color_data = 12'b001110100111;
		16'b0110111011001100: color_data = 12'b001110100111;
		16'b0110111011001101: color_data = 12'b001110100111;
		16'b0110111011001110: color_data = 12'b001110100111;
		16'b0110111011001111: color_data = 12'b001110100111;
		16'b0110111011010000: color_data = 12'b001110100111;
		16'b0110111011010001: color_data = 12'b001110100111;
		16'b0110111011010010: color_data = 12'b001110100111;
		16'b0110111011010011: color_data = 12'b001110100111;
		16'b0110111011010100: color_data = 12'b001110100111;
		16'b0110111011010101: color_data = 12'b001110100111;
		16'b0110111011010110: color_data = 12'b001110100111;
		16'b0110111011010111: color_data = 12'b001110100111;
		16'b0110111011011000: color_data = 12'b001110100111;
		16'b0110111011011001: color_data = 12'b001110100111;
		16'b0110111011011010: color_data = 12'b001110100111;
		16'b0110111011011011: color_data = 12'b001110100111;
		16'b0110111011011100: color_data = 12'b001110100111;
		16'b0110111011011101: color_data = 12'b001110100111;
		16'b0110111011011110: color_data = 12'b001110100111;
		16'b0110111011011111: color_data = 12'b001110100111;
		16'b0110111011100000: color_data = 12'b001110100111;
		16'b0110111011100001: color_data = 12'b001110100111;
		16'b0110111011100010: color_data = 12'b001110100111;
		16'b0110111011110110: color_data = 12'b001110100111;
		16'b0110111011110111: color_data = 12'b001110100111;
		16'b0110111011111000: color_data = 12'b001110100111;
		16'b0110111011111001: color_data = 12'b001110100111;
		16'b0110111011111010: color_data = 12'b001110100111;
		16'b0110111011111011: color_data = 12'b001110100111;
		16'b0110111011111100: color_data = 12'b001110100111;
		16'b0110111011111101: color_data = 12'b001110100111;
		16'b0110111011111110: color_data = 12'b001110100111;
		16'b0110111011111111: color_data = 12'b001110100111;
		16'b0110111100000000: color_data = 12'b001110100111;
		16'b0110111100000001: color_data = 12'b001110100111;
		16'b0110111100011010: color_data = 12'b001110100111;
		16'b0110111100011011: color_data = 12'b001110100111;
		16'b0110111100011100: color_data = 12'b001110100111;
		16'b0110111100011101: color_data = 12'b001110100111;
		16'b0110111100011110: color_data = 12'b001110100111;
		16'b0110111100011111: color_data = 12'b001110100111;
		16'b0110111100100000: color_data = 12'b001110100111;
		16'b0110111100100001: color_data = 12'b001110100111;
		16'b0110111100100010: color_data = 12'b001110100111;
		16'b0110111100100011: color_data = 12'b001110100111;
		16'b0110111100100100: color_data = 12'b001110100111;
		16'b0110111100100101: color_data = 12'b001110100111;
		16'b0110111100100110: color_data = 12'b001110100111;
		16'b0110111100101101: color_data = 12'b001110100111;
		16'b0110111100101110: color_data = 12'b001110100111;
		16'b0110111100101111: color_data = 12'b001110100111;
		16'b0110111100110000: color_data = 12'b001110100111;
		16'b0110111100110001: color_data = 12'b001110100111;
		16'b0110111100110010: color_data = 12'b001110100111;
		16'b0110111100110011: color_data = 12'b001110100111;
		16'b0110111100110100: color_data = 12'b001110100111;
		16'b0110111100110101: color_data = 12'b001110100111;
		16'b0110111100110110: color_data = 12'b001110100111;
		16'b0110111100110111: color_data = 12'b001110100111;
		16'b0110111100111000: color_data = 12'b001110100111;
		16'b0110111101000101: color_data = 12'b001110100111;
		16'b0110111101000110: color_data = 12'b001110100111;
		16'b0110111101000111: color_data = 12'b001110100111;
		16'b0110111101001000: color_data = 12'b001110100111;
		16'b0110111101001001: color_data = 12'b001110100111;
		16'b0110111101001010: color_data = 12'b001110100111;
		16'b0110111101001011: color_data = 12'b001110100111;
		16'b0110111101001100: color_data = 12'b001110100111;
		16'b0110111101001101: color_data = 12'b001110100111;
		16'b0110111101001110: color_data = 12'b001110100111;
		16'b0110111101001111: color_data = 12'b001110100111;
		16'b0110111101010000: color_data = 12'b001110100111;
		16'b0110111101010001: color_data = 12'b001110100111;
		16'b0110111101011000: color_data = 12'b001110100111;
		16'b0110111101011001: color_data = 12'b001110100111;
		16'b0110111101011010: color_data = 12'b001110100111;
		16'b0110111101011011: color_data = 12'b001110100111;
		16'b0110111101011100: color_data = 12'b001110100111;
		16'b0110111101011101: color_data = 12'b001110100111;
		16'b0110111101011110: color_data = 12'b001110100111;
		16'b0110111101011111: color_data = 12'b001110100111;
		16'b0110111101100000: color_data = 12'b001110100111;
		16'b0110111101100001: color_data = 12'b001110100111;
		16'b0110111101100010: color_data = 12'b001110100111;
		16'b0110111101100011: color_data = 12'b001110100111;
		16'b0110111101110000: color_data = 12'b001110100111;
		16'b0110111101110001: color_data = 12'b001110100111;
		16'b0110111101110010: color_data = 12'b001110100111;
		16'b0110111101110011: color_data = 12'b001110100111;
		16'b0110111101110100: color_data = 12'b001110100111;
		16'b0110111101110101: color_data = 12'b001110100111;
		16'b0110111101110110: color_data = 12'b001110100111;
		16'b0110111101110111: color_data = 12'b001110100111;
		16'b0110111101111000: color_data = 12'b001110100111;
		16'b0110111101111001: color_data = 12'b001110100111;
		16'b0110111101111010: color_data = 12'b001110100111;
		16'b0110111101111011: color_data = 12'b001110100111;
		16'b0111000000000000: color_data = 12'b001110100111;
		16'b0111000000000001: color_data = 12'b001110100111;
		16'b0111000000000010: color_data = 12'b001110100111;
		16'b0111000000000011: color_data = 12'b001110100111;
		16'b0111000000000100: color_data = 12'b001110100111;
		16'b0111000000000101: color_data = 12'b001110100111;
		16'b0111000000000110: color_data = 12'b001110100111;
		16'b0111000000000111: color_data = 12'b001110100111;
		16'b0111000000001000: color_data = 12'b001110100111;
		16'b0111000000001001: color_data = 12'b001110100111;
		16'b0111000000001010: color_data = 12'b001110100111;
		16'b0111000000001011: color_data = 12'b001110100111;
		16'b0111000000001100: color_data = 12'b001110100111;
		16'b0111000000101011: color_data = 12'b001110100111;
		16'b0111000000101100: color_data = 12'b001110100111;
		16'b0111000000101101: color_data = 12'b001110100111;
		16'b0111000000101110: color_data = 12'b001110100111;
		16'b0111000000101111: color_data = 12'b001110100111;
		16'b0111000000110000: color_data = 12'b001110100111;
		16'b0111000000110001: color_data = 12'b001110100111;
		16'b0111000000110010: color_data = 12'b001110100111;
		16'b0111000000110011: color_data = 12'b001110100111;
		16'b0111000000110100: color_data = 12'b001110100111;
		16'b0111000000110101: color_data = 12'b001110100111;
		16'b0111000000110110: color_data = 12'b001110100111;
		16'b0111000000110111: color_data = 12'b001110100111;
		16'b0111000000111000: color_data = 12'b001110100111;
		16'b0111000000111001: color_data = 12'b001110100111;
		16'b0111000000111010: color_data = 12'b001110100111;
		16'b0111000000111011: color_data = 12'b001110100111;
		16'b0111000000111100: color_data = 12'b001110100111;
		16'b0111000000111101: color_data = 12'b001110100111;
		16'b0111000000111110: color_data = 12'b001110100111;
		16'b0111000000111111: color_data = 12'b001110100111;
		16'b0111000001000000: color_data = 12'b001110100111;
		16'b0111000001000001: color_data = 12'b001110100111;
		16'b0111000001000010: color_data = 12'b001110100111;
		16'b0111000001000011: color_data = 12'b001110100111;
		16'b0111000001000100: color_data = 12'b001110100111;
		16'b0111000001000101: color_data = 12'b001110100111;
		16'b0111000001000110: color_data = 12'b001110100111;
		16'b0111000001000111: color_data = 12'b001110100111;
		16'b0111000001001000: color_data = 12'b001110100111;
		16'b0111000001001001: color_data = 12'b001110100111;
		16'b0111000001001010: color_data = 12'b001110100111;
		16'b0111000001001011: color_data = 12'b001110100111;
		16'b0111000001001100: color_data = 12'b001110100111;
		16'b0111000001001101: color_data = 12'b001110100111;
		16'b0111000001001110: color_data = 12'b001110100111;
		16'b0111000001001111: color_data = 12'b001110100111;
		16'b0111000001011100: color_data = 12'b001110100111;
		16'b0111000001011101: color_data = 12'b001110100111;
		16'b0111000001011110: color_data = 12'b001110100111;
		16'b0111000001011111: color_data = 12'b001110100111;
		16'b0111000001100000: color_data = 12'b001110100111;
		16'b0111000001100001: color_data = 12'b001110100111;
		16'b0111000001100010: color_data = 12'b001110100111;
		16'b0111000001100011: color_data = 12'b001110100111;
		16'b0111000001100100: color_data = 12'b001110100111;
		16'b0111000001100101: color_data = 12'b001110100111;
		16'b0111000001100110: color_data = 12'b001110100111;
		16'b0111000001100111: color_data = 12'b001110100111;
		16'b0111000001101000: color_data = 12'b001110100111;
		16'b0111000001110101: color_data = 12'b001110100111;
		16'b0111000001110110: color_data = 12'b001110100111;
		16'b0111000001110111: color_data = 12'b001110100111;
		16'b0111000001111000: color_data = 12'b001110100111;
		16'b0111000001111001: color_data = 12'b001110100111;
		16'b0111000001111010: color_data = 12'b001110100111;
		16'b0111000001111011: color_data = 12'b001110100111;
		16'b0111000001111100: color_data = 12'b001110100111;
		16'b0111000001111101: color_data = 12'b001110100111;
		16'b0111000001111110: color_data = 12'b001110100111;
		16'b0111000001111111: color_data = 12'b001110100111;
		16'b0111000010000000: color_data = 12'b001110100111;
		16'b0111000010001101: color_data = 12'b001110100111;
		16'b0111000010001110: color_data = 12'b001110100111;
		16'b0111000010001111: color_data = 12'b001110100111;
		16'b0111000010010000: color_data = 12'b001110100111;
		16'b0111000010010001: color_data = 12'b001110100111;
		16'b0111000010010010: color_data = 12'b001110100111;
		16'b0111000010010011: color_data = 12'b001110100111;
		16'b0111000010010100: color_data = 12'b001110100111;
		16'b0111000010010101: color_data = 12'b001110100111;
		16'b0111000010010110: color_data = 12'b001110100111;
		16'b0111000010010111: color_data = 12'b001110100111;
		16'b0111000010011000: color_data = 12'b001110100111;
		16'b0111000010011001: color_data = 12'b001110100111;
		16'b0111000010100000: color_data = 12'b001110100111;
		16'b0111000010100001: color_data = 12'b001110100111;
		16'b0111000010100010: color_data = 12'b001110100111;
		16'b0111000010100011: color_data = 12'b001110100111;
		16'b0111000010100100: color_data = 12'b001110100111;
		16'b0111000010100101: color_data = 12'b001110100111;
		16'b0111000010100110: color_data = 12'b001110100111;
		16'b0111000010100111: color_data = 12'b001110100111;
		16'b0111000010101000: color_data = 12'b001110100111;
		16'b0111000010101001: color_data = 12'b001110100111;
		16'b0111000010101010: color_data = 12'b001110100111;
		16'b0111000010101011: color_data = 12'b001110100111;
		16'b0111000010111000: color_data = 12'b001110100111;
		16'b0111000010111001: color_data = 12'b001110100111;
		16'b0111000010111010: color_data = 12'b001110100111;
		16'b0111000010111011: color_data = 12'b001110100111;
		16'b0111000010111100: color_data = 12'b001110100111;
		16'b0111000010111101: color_data = 12'b001110100111;
		16'b0111000010111110: color_data = 12'b001110100111;
		16'b0111000010111111: color_data = 12'b001110100111;
		16'b0111000011000000: color_data = 12'b001110100111;
		16'b0111000011000001: color_data = 12'b001110100111;
		16'b0111000011000010: color_data = 12'b001110100111;
		16'b0111000011000011: color_data = 12'b001110100111;
		16'b0111000011000100: color_data = 12'b001110100111;
		16'b0111000011001011: color_data = 12'b001110100111;
		16'b0111000011001100: color_data = 12'b001110100111;
		16'b0111000011001101: color_data = 12'b001110100111;
		16'b0111000011001110: color_data = 12'b001110100111;
		16'b0111000011001111: color_data = 12'b001110100111;
		16'b0111000011010000: color_data = 12'b001110100111;
		16'b0111000011010001: color_data = 12'b001110100111;
		16'b0111000011010010: color_data = 12'b001110100111;
		16'b0111000011010011: color_data = 12'b001110100111;
		16'b0111000011010100: color_data = 12'b001110100111;
		16'b0111000011010101: color_data = 12'b001110100111;
		16'b0111000011010110: color_data = 12'b001110100111;
		16'b0111000011010111: color_data = 12'b001110100111;
		16'b0111000011011000: color_data = 12'b001110100111;
		16'b0111000011011001: color_data = 12'b001110100111;
		16'b0111000011011010: color_data = 12'b001110100111;
		16'b0111000011011011: color_data = 12'b001110100111;
		16'b0111000011011100: color_data = 12'b001110100111;
		16'b0111000011011101: color_data = 12'b001110100111;
		16'b0111000011011110: color_data = 12'b001110100111;
		16'b0111000011011111: color_data = 12'b001110100111;
		16'b0111000011100000: color_data = 12'b001110100111;
		16'b0111000011100001: color_data = 12'b001110100111;
		16'b0111000011100010: color_data = 12'b001110100111;
		16'b0111000011110110: color_data = 12'b001110100111;
		16'b0111000011110111: color_data = 12'b001110100111;
		16'b0111000011111000: color_data = 12'b001110100111;
		16'b0111000011111001: color_data = 12'b001110100111;
		16'b0111000011111010: color_data = 12'b001110100111;
		16'b0111000011111011: color_data = 12'b001110100111;
		16'b0111000011111100: color_data = 12'b001110100111;
		16'b0111000011111101: color_data = 12'b001110100111;
		16'b0111000011111110: color_data = 12'b001110100111;
		16'b0111000011111111: color_data = 12'b001110100111;
		16'b0111000100000000: color_data = 12'b001110100111;
		16'b0111000100000001: color_data = 12'b001110100111;
		16'b0111000100011010: color_data = 12'b001110100111;
		16'b0111000100011011: color_data = 12'b001110100111;
		16'b0111000100011100: color_data = 12'b001110100111;
		16'b0111000100011101: color_data = 12'b001110100111;
		16'b0111000100011110: color_data = 12'b001110100111;
		16'b0111000100011111: color_data = 12'b001110100111;
		16'b0111000100100000: color_data = 12'b001110100111;
		16'b0111000100100001: color_data = 12'b001110100111;
		16'b0111000100100010: color_data = 12'b001110100111;
		16'b0111000100100011: color_data = 12'b001110100111;
		16'b0111000100100100: color_data = 12'b001110100111;
		16'b0111000100100101: color_data = 12'b001110100111;
		16'b0111000100100110: color_data = 12'b001110100111;
		16'b0111000100101101: color_data = 12'b001110100111;
		16'b0111000100101110: color_data = 12'b001110100111;
		16'b0111000100101111: color_data = 12'b001110100111;
		16'b0111000100110000: color_data = 12'b001110100111;
		16'b0111000100110001: color_data = 12'b001110100111;
		16'b0111000100110010: color_data = 12'b001110100111;
		16'b0111000100110011: color_data = 12'b001110100111;
		16'b0111000100110100: color_data = 12'b001110100111;
		16'b0111000100110101: color_data = 12'b001110100111;
		16'b0111000100110110: color_data = 12'b001110100111;
		16'b0111000100110111: color_data = 12'b001110100111;
		16'b0111000100111000: color_data = 12'b001110100111;
		16'b0111000101000101: color_data = 12'b001110100111;
		16'b0111000101000110: color_data = 12'b001110100111;
		16'b0111000101000111: color_data = 12'b001110100111;
		16'b0111000101001000: color_data = 12'b001110100111;
		16'b0111000101001001: color_data = 12'b001110100111;
		16'b0111000101001010: color_data = 12'b001110100111;
		16'b0111000101001011: color_data = 12'b001110100111;
		16'b0111000101001100: color_data = 12'b001110100111;
		16'b0111000101001101: color_data = 12'b001110100111;
		16'b0111000101001110: color_data = 12'b001110100111;
		16'b0111000101001111: color_data = 12'b001110100111;
		16'b0111000101010000: color_data = 12'b001110100111;
		16'b0111000101010001: color_data = 12'b001110100111;
		16'b0111000101011000: color_data = 12'b001110100111;
		16'b0111000101011001: color_data = 12'b001110100111;
		16'b0111000101011010: color_data = 12'b001110100111;
		16'b0111000101011011: color_data = 12'b001110100111;
		16'b0111000101011100: color_data = 12'b001110100111;
		16'b0111000101011101: color_data = 12'b001110100111;
		16'b0111000101011110: color_data = 12'b001110100111;
		16'b0111000101011111: color_data = 12'b001110100111;
		16'b0111000101100000: color_data = 12'b001110100111;
		16'b0111000101100001: color_data = 12'b001110100111;
		16'b0111000101100010: color_data = 12'b001110100111;
		16'b0111000101100011: color_data = 12'b001110100111;
		16'b0111000101110000: color_data = 12'b001110100111;
		16'b0111000101110001: color_data = 12'b001110100111;
		16'b0111000101110010: color_data = 12'b001110100111;
		16'b0111000101110011: color_data = 12'b001110100111;
		16'b0111000101110100: color_data = 12'b001110100111;
		16'b0111000101110101: color_data = 12'b001110100111;
		16'b0111000101110110: color_data = 12'b001110100111;
		16'b0111000101110111: color_data = 12'b001110100111;
		16'b0111000101111000: color_data = 12'b001110100111;
		16'b0111000101111001: color_data = 12'b001110100111;
		16'b0111000101111010: color_data = 12'b001110100111;
		16'b0111000101111011: color_data = 12'b001110100111;
		16'b0111001000000000: color_data = 12'b001110100111;
		16'b0111001000000001: color_data = 12'b001110100111;
		16'b0111001000000010: color_data = 12'b001110100111;
		16'b0111001000000011: color_data = 12'b001110100111;
		16'b0111001000000100: color_data = 12'b001110100111;
		16'b0111001000000101: color_data = 12'b001110100111;
		16'b0111001000000110: color_data = 12'b001110100111;
		16'b0111001000000111: color_data = 12'b001110100111;
		16'b0111001000001000: color_data = 12'b001110100111;
		16'b0111001000001001: color_data = 12'b001110100111;
		16'b0111001000001010: color_data = 12'b001110100111;
		16'b0111001000001011: color_data = 12'b001110100111;
		16'b0111001000001100: color_data = 12'b001110100111;
		16'b0111001000101011: color_data = 12'b001110100111;
		16'b0111001000101100: color_data = 12'b001110100111;
		16'b0111001000101101: color_data = 12'b001110100111;
		16'b0111001000101110: color_data = 12'b001110100111;
		16'b0111001000101111: color_data = 12'b001110100111;
		16'b0111001000110000: color_data = 12'b001110100111;
		16'b0111001000110001: color_data = 12'b001110100111;
		16'b0111001000110010: color_data = 12'b001110100111;
		16'b0111001000110011: color_data = 12'b001110100111;
		16'b0111001000110100: color_data = 12'b001110100111;
		16'b0111001000110101: color_data = 12'b001110100111;
		16'b0111001000110110: color_data = 12'b001110100111;
		16'b0111001000110111: color_data = 12'b001110100111;
		16'b0111001000111000: color_data = 12'b001110100111;
		16'b0111001000111001: color_data = 12'b001110100111;
		16'b0111001000111010: color_data = 12'b001110100111;
		16'b0111001000111011: color_data = 12'b001110100111;
		16'b0111001000111100: color_data = 12'b001110100111;
		16'b0111001000111101: color_data = 12'b001110100111;
		16'b0111001000111110: color_data = 12'b001110100111;
		16'b0111001000111111: color_data = 12'b001110100111;
		16'b0111001001000000: color_data = 12'b001110100111;
		16'b0111001001000001: color_data = 12'b001110100111;
		16'b0111001001000010: color_data = 12'b001110100111;
		16'b0111001001000011: color_data = 12'b001110100111;
		16'b0111001001000100: color_data = 12'b001110100111;
		16'b0111001001000101: color_data = 12'b001110100111;
		16'b0111001001000110: color_data = 12'b001110100111;
		16'b0111001001000111: color_data = 12'b001110100111;
		16'b0111001001001000: color_data = 12'b001110100111;
		16'b0111001001001001: color_data = 12'b001110100111;
		16'b0111001001001010: color_data = 12'b001110100111;
		16'b0111001001001011: color_data = 12'b001110100111;
		16'b0111001001001100: color_data = 12'b001110100111;
		16'b0111001001001101: color_data = 12'b001110100111;
		16'b0111001001001110: color_data = 12'b001110100111;
		16'b0111001001001111: color_data = 12'b001110100111;
		16'b0111001001011100: color_data = 12'b001110100111;
		16'b0111001001011101: color_data = 12'b001110100111;
		16'b0111001001011110: color_data = 12'b001110100111;
		16'b0111001001011111: color_data = 12'b001110100111;
		16'b0111001001100000: color_data = 12'b001110100111;
		16'b0111001001100001: color_data = 12'b001110100111;
		16'b0111001001100010: color_data = 12'b001110100111;
		16'b0111001001100011: color_data = 12'b001110100111;
		16'b0111001001100100: color_data = 12'b001110100111;
		16'b0111001001100101: color_data = 12'b001110100111;
		16'b0111001001100110: color_data = 12'b001110100111;
		16'b0111001001100111: color_data = 12'b001110100111;
		16'b0111001001101000: color_data = 12'b001110100111;
		16'b0111001001110101: color_data = 12'b001110100111;
		16'b0111001001110110: color_data = 12'b001110100111;
		16'b0111001001110111: color_data = 12'b001110100111;
		16'b0111001001111000: color_data = 12'b001110100111;
		16'b0111001001111001: color_data = 12'b001110100111;
		16'b0111001001111010: color_data = 12'b001110100111;
		16'b0111001001111011: color_data = 12'b001110100111;
		16'b0111001001111100: color_data = 12'b001110100111;
		16'b0111001001111101: color_data = 12'b001110100111;
		16'b0111001001111110: color_data = 12'b001110100111;
		16'b0111001001111111: color_data = 12'b001110100111;
		16'b0111001010000000: color_data = 12'b001110100111;
		16'b0111001010001101: color_data = 12'b001110100111;
		16'b0111001010001110: color_data = 12'b001110100111;
		16'b0111001010001111: color_data = 12'b001110100111;
		16'b0111001010010000: color_data = 12'b001110100111;
		16'b0111001010010001: color_data = 12'b001110100111;
		16'b0111001010010010: color_data = 12'b001110100111;
		16'b0111001010010011: color_data = 12'b001110100111;
		16'b0111001010010100: color_data = 12'b001110100111;
		16'b0111001010010101: color_data = 12'b001110100111;
		16'b0111001010010110: color_data = 12'b001110100111;
		16'b0111001010010111: color_data = 12'b001110100111;
		16'b0111001010011000: color_data = 12'b001110100111;
		16'b0111001010011001: color_data = 12'b001110100111;
		16'b0111001010100000: color_data = 12'b001110100111;
		16'b0111001010100001: color_data = 12'b001110100111;
		16'b0111001010100010: color_data = 12'b001110100111;
		16'b0111001010100011: color_data = 12'b001110100111;
		16'b0111001010100100: color_data = 12'b001110100111;
		16'b0111001010100101: color_data = 12'b001110100111;
		16'b0111001010100110: color_data = 12'b001110100111;
		16'b0111001010100111: color_data = 12'b001110100111;
		16'b0111001010101000: color_data = 12'b001110100111;
		16'b0111001010101001: color_data = 12'b001110100111;
		16'b0111001010101010: color_data = 12'b001110100111;
		16'b0111001010101011: color_data = 12'b001110100111;
		16'b0111001010111000: color_data = 12'b001110100111;
		16'b0111001010111001: color_data = 12'b001110100111;
		16'b0111001010111010: color_data = 12'b001110100111;
		16'b0111001010111011: color_data = 12'b001110100111;
		16'b0111001010111100: color_data = 12'b001110100111;
		16'b0111001010111101: color_data = 12'b001110100111;
		16'b0111001010111110: color_data = 12'b001110100111;
		16'b0111001010111111: color_data = 12'b001110100111;
		16'b0111001011000000: color_data = 12'b001110100111;
		16'b0111001011000001: color_data = 12'b001110100111;
		16'b0111001011000010: color_data = 12'b001110100111;
		16'b0111001011000011: color_data = 12'b001110100111;
		16'b0111001011000100: color_data = 12'b001110100111;
		16'b0111001011001011: color_data = 12'b001110100111;
		16'b0111001011001100: color_data = 12'b001110100111;
		16'b0111001011001101: color_data = 12'b001110100111;
		16'b0111001011001110: color_data = 12'b001110100111;
		16'b0111001011001111: color_data = 12'b001110100111;
		16'b0111001011010000: color_data = 12'b001110100111;
		16'b0111001011010001: color_data = 12'b001110100111;
		16'b0111001011010010: color_data = 12'b001110100111;
		16'b0111001011010011: color_data = 12'b001110100111;
		16'b0111001011010100: color_data = 12'b001110100111;
		16'b0111001011010101: color_data = 12'b001110100111;
		16'b0111001011010110: color_data = 12'b001110100111;
		16'b0111001011010111: color_data = 12'b001110100111;
		16'b0111001011011000: color_data = 12'b001110100111;
		16'b0111001011011001: color_data = 12'b001110100111;
		16'b0111001011011010: color_data = 12'b001110100111;
		16'b0111001011011011: color_data = 12'b001110100111;
		16'b0111001011011100: color_data = 12'b001110100111;
		16'b0111001011011101: color_data = 12'b001110100111;
		16'b0111001011011110: color_data = 12'b001110100111;
		16'b0111001011011111: color_data = 12'b001110100111;
		16'b0111001011100000: color_data = 12'b001110100111;
		16'b0111001011100001: color_data = 12'b001110100111;
		16'b0111001011100010: color_data = 12'b001110100111;
		16'b0111001011110110: color_data = 12'b001110100111;
		16'b0111001011110111: color_data = 12'b001110100111;
		16'b0111001011111000: color_data = 12'b001110100111;
		16'b0111001011111001: color_data = 12'b001110100111;
		16'b0111001011111010: color_data = 12'b001110100111;
		16'b0111001011111011: color_data = 12'b001110100111;
		16'b0111001011111100: color_data = 12'b001110100111;
		16'b0111001011111101: color_data = 12'b001110100111;
		16'b0111001011111110: color_data = 12'b001110100111;
		16'b0111001011111111: color_data = 12'b001110100111;
		16'b0111001100000000: color_data = 12'b001110100111;
		16'b0111001100000001: color_data = 12'b001110100111;
		16'b0111001100011010: color_data = 12'b001110100111;
		16'b0111001100011011: color_data = 12'b001110100111;
		16'b0111001100011100: color_data = 12'b001110100111;
		16'b0111001100011101: color_data = 12'b001110100111;
		16'b0111001100011110: color_data = 12'b001110100111;
		16'b0111001100011111: color_data = 12'b001110100111;
		16'b0111001100100000: color_data = 12'b001110100111;
		16'b0111001100100001: color_data = 12'b001110100111;
		16'b0111001100100010: color_data = 12'b001110100111;
		16'b0111001100100011: color_data = 12'b001110100111;
		16'b0111001100100100: color_data = 12'b001110100111;
		16'b0111001100100101: color_data = 12'b001110100111;
		16'b0111001100100110: color_data = 12'b001110100111;
		16'b0111001100101101: color_data = 12'b001110100111;
		16'b0111001100101110: color_data = 12'b001110100111;
		16'b0111001100101111: color_data = 12'b001110100111;
		16'b0111001100110000: color_data = 12'b001110100111;
		16'b0111001100110001: color_data = 12'b001110100111;
		16'b0111001100110010: color_data = 12'b001110100111;
		16'b0111001100110011: color_data = 12'b001110100111;
		16'b0111001100110100: color_data = 12'b001110100111;
		16'b0111001100110101: color_data = 12'b001110100111;
		16'b0111001100110110: color_data = 12'b001110100111;
		16'b0111001100110111: color_data = 12'b001110100111;
		16'b0111001100111000: color_data = 12'b001110100111;
		16'b0111001101000101: color_data = 12'b001110100111;
		16'b0111001101000110: color_data = 12'b001110100111;
		16'b0111001101000111: color_data = 12'b001110100111;
		16'b0111001101001000: color_data = 12'b001110100111;
		16'b0111001101001001: color_data = 12'b001110100111;
		16'b0111001101001010: color_data = 12'b001110100111;
		16'b0111001101001011: color_data = 12'b001110100111;
		16'b0111001101001100: color_data = 12'b001110100111;
		16'b0111001101001101: color_data = 12'b001110100111;
		16'b0111001101001110: color_data = 12'b001110100111;
		16'b0111001101001111: color_data = 12'b001110100111;
		16'b0111001101010000: color_data = 12'b001110100111;
		16'b0111001101010001: color_data = 12'b001110100111;
		16'b0111001101011000: color_data = 12'b001110100111;
		16'b0111001101011001: color_data = 12'b001110100111;
		16'b0111001101011010: color_data = 12'b001110100111;
		16'b0111001101011011: color_data = 12'b001110100111;
		16'b0111001101011100: color_data = 12'b001110100111;
		16'b0111001101011101: color_data = 12'b001110100111;
		16'b0111001101011110: color_data = 12'b001110100111;
		16'b0111001101011111: color_data = 12'b001110100111;
		16'b0111001101100000: color_data = 12'b001110100111;
		16'b0111001101100001: color_data = 12'b001110100111;
		16'b0111001101100010: color_data = 12'b001110100111;
		16'b0111001101100011: color_data = 12'b001110100111;
		16'b0111001101110000: color_data = 12'b001110100111;
		16'b0111001101110001: color_data = 12'b001110100111;
		16'b0111001101110010: color_data = 12'b001110100111;
		16'b0111001101110011: color_data = 12'b001110100111;
		16'b0111001101110100: color_data = 12'b001110100111;
		16'b0111001101110101: color_data = 12'b001110100111;
		16'b0111001101110110: color_data = 12'b001110100111;
		16'b0111001101110111: color_data = 12'b001110100111;
		16'b0111001101111000: color_data = 12'b001110100111;
		16'b0111001101111001: color_data = 12'b001110100111;
		16'b0111001101111010: color_data = 12'b001110100111;
		16'b0111001101111011: color_data = 12'b001110100111;
		16'b0111010000000000: color_data = 12'b001110100111;
		16'b0111010000000001: color_data = 12'b001110100111;
		16'b0111010000000010: color_data = 12'b001110100111;
		16'b0111010000000011: color_data = 12'b001110100111;
		16'b0111010000000100: color_data = 12'b001110100111;
		16'b0111010000000101: color_data = 12'b001110100111;
		16'b0111010000000110: color_data = 12'b001110100111;
		16'b0111010000000111: color_data = 12'b001110100111;
		16'b0111010000001000: color_data = 12'b001110100111;
		16'b0111010000001001: color_data = 12'b001110100111;
		16'b0111010000001010: color_data = 12'b001110100111;
		16'b0111010000001011: color_data = 12'b001110100111;
		16'b0111010000001100: color_data = 12'b001110100111;
		16'b0111010000101011: color_data = 12'b001110100111;
		16'b0111010000101100: color_data = 12'b001110100111;
		16'b0111010000101101: color_data = 12'b001110100111;
		16'b0111010000101110: color_data = 12'b001110100111;
		16'b0111010000101111: color_data = 12'b001110100111;
		16'b0111010000110000: color_data = 12'b001110100111;
		16'b0111010000110001: color_data = 12'b001110100111;
		16'b0111010000110010: color_data = 12'b001110100111;
		16'b0111010000110011: color_data = 12'b001110100111;
		16'b0111010000110100: color_data = 12'b001110100111;
		16'b0111010000110101: color_data = 12'b001110100111;
		16'b0111010000110110: color_data = 12'b001110100111;
		16'b0111010000110111: color_data = 12'b001110100111;
		16'b0111010000111000: color_data = 12'b001110100111;
		16'b0111010000111001: color_data = 12'b001110100111;
		16'b0111010000111010: color_data = 12'b001110100111;
		16'b0111010000111011: color_data = 12'b001110100111;
		16'b0111010000111100: color_data = 12'b001110100111;
		16'b0111010000111101: color_data = 12'b001110100111;
		16'b0111010000111110: color_data = 12'b001110100111;
		16'b0111010000111111: color_data = 12'b001110100111;
		16'b0111010001000000: color_data = 12'b001110100111;
		16'b0111010001000001: color_data = 12'b001110100111;
		16'b0111010001000010: color_data = 12'b001110100111;
		16'b0111010001000011: color_data = 12'b001110100111;
		16'b0111010001000100: color_data = 12'b001110100111;
		16'b0111010001000101: color_data = 12'b001110100111;
		16'b0111010001000110: color_data = 12'b001110100111;
		16'b0111010001000111: color_data = 12'b001110100111;
		16'b0111010001001000: color_data = 12'b001110100111;
		16'b0111010001001001: color_data = 12'b001110100111;
		16'b0111010001001010: color_data = 12'b001110100111;
		16'b0111010001001011: color_data = 12'b001110100111;
		16'b0111010001001100: color_data = 12'b001110100111;
		16'b0111010001001101: color_data = 12'b001110100111;
		16'b0111010001001110: color_data = 12'b001110100111;
		16'b0111010001001111: color_data = 12'b001110100111;
		16'b0111010001011100: color_data = 12'b001110100111;
		16'b0111010001011101: color_data = 12'b001110100111;
		16'b0111010001011110: color_data = 12'b001110100111;
		16'b0111010001011111: color_data = 12'b001110100111;
		16'b0111010001100000: color_data = 12'b001110100111;
		16'b0111010001100001: color_data = 12'b001110100111;
		16'b0111010001100010: color_data = 12'b001110100111;
		16'b0111010001100011: color_data = 12'b001110100111;
		16'b0111010001100100: color_data = 12'b001110100111;
		16'b0111010001100101: color_data = 12'b001110100111;
		16'b0111010001100110: color_data = 12'b001110100111;
		16'b0111010001100111: color_data = 12'b001110100111;
		16'b0111010001101000: color_data = 12'b001110100111;
		16'b0111010001110101: color_data = 12'b001110100111;
		16'b0111010001110110: color_data = 12'b001110100111;
		16'b0111010001110111: color_data = 12'b001110100111;
		16'b0111010001111000: color_data = 12'b001110100111;
		16'b0111010001111001: color_data = 12'b001110100111;
		16'b0111010001111010: color_data = 12'b001110100111;
		16'b0111010001111011: color_data = 12'b001110100111;
		16'b0111010001111100: color_data = 12'b001110100111;
		16'b0111010001111101: color_data = 12'b001110100111;
		16'b0111010001111110: color_data = 12'b001110100111;
		16'b0111010001111111: color_data = 12'b001110100111;
		16'b0111010010000000: color_data = 12'b001110100111;
		16'b0111010010001101: color_data = 12'b001110100111;
		16'b0111010010001110: color_data = 12'b001110100111;
		16'b0111010010001111: color_data = 12'b001110100111;
		16'b0111010010010000: color_data = 12'b001110100111;
		16'b0111010010010001: color_data = 12'b001110100111;
		16'b0111010010010010: color_data = 12'b001110100111;
		16'b0111010010010011: color_data = 12'b001110100111;
		16'b0111010010010100: color_data = 12'b001110100111;
		16'b0111010010010101: color_data = 12'b001110100111;
		16'b0111010010010110: color_data = 12'b001110100111;
		16'b0111010010010111: color_data = 12'b001110100111;
		16'b0111010010011000: color_data = 12'b001110100111;
		16'b0111010010011001: color_data = 12'b001110100111;
		16'b0111010010100000: color_data = 12'b001110100111;
		16'b0111010010100001: color_data = 12'b001110100111;
		16'b0111010010100010: color_data = 12'b001110100111;
		16'b0111010010100011: color_data = 12'b001110100111;
		16'b0111010010100100: color_data = 12'b001110100111;
		16'b0111010010100101: color_data = 12'b001110100111;
		16'b0111010010100110: color_data = 12'b001110100111;
		16'b0111010010100111: color_data = 12'b001110100111;
		16'b0111010010101000: color_data = 12'b001110100111;
		16'b0111010010101001: color_data = 12'b001110100111;
		16'b0111010010101010: color_data = 12'b001110100111;
		16'b0111010010101011: color_data = 12'b001110100111;
		16'b0111010010111000: color_data = 12'b001110100111;
		16'b0111010010111001: color_data = 12'b001110100111;
		16'b0111010010111010: color_data = 12'b001110100111;
		16'b0111010010111011: color_data = 12'b001110100111;
		16'b0111010010111100: color_data = 12'b001110100111;
		16'b0111010010111101: color_data = 12'b001110100111;
		16'b0111010010111110: color_data = 12'b001110100111;
		16'b0111010010111111: color_data = 12'b001110100111;
		16'b0111010011000000: color_data = 12'b001110100111;
		16'b0111010011000001: color_data = 12'b001110100111;
		16'b0111010011000010: color_data = 12'b001110100111;
		16'b0111010011000011: color_data = 12'b001110100111;
		16'b0111010011000100: color_data = 12'b001110100111;
		16'b0111010011001011: color_data = 12'b001110100111;
		16'b0111010011001100: color_data = 12'b001110100111;
		16'b0111010011001101: color_data = 12'b001110100111;
		16'b0111010011001110: color_data = 12'b001110100111;
		16'b0111010011001111: color_data = 12'b001110100111;
		16'b0111010011010000: color_data = 12'b001110100111;
		16'b0111010011010001: color_data = 12'b001110100111;
		16'b0111010011010010: color_data = 12'b001110100111;
		16'b0111010011010011: color_data = 12'b001110100111;
		16'b0111010011010100: color_data = 12'b001110100111;
		16'b0111010011010101: color_data = 12'b001110100111;
		16'b0111010011010110: color_data = 12'b001110100111;
		16'b0111010011010111: color_data = 12'b001110100111;
		16'b0111010011011000: color_data = 12'b001110100111;
		16'b0111010011011001: color_data = 12'b001110100111;
		16'b0111010011011010: color_data = 12'b001110100111;
		16'b0111010011011011: color_data = 12'b001110100111;
		16'b0111010011011100: color_data = 12'b001110100111;
		16'b0111010011011101: color_data = 12'b001110100111;
		16'b0111010011011110: color_data = 12'b001110100111;
		16'b0111010011011111: color_data = 12'b001110100111;
		16'b0111010011100000: color_data = 12'b001110100111;
		16'b0111010011100001: color_data = 12'b001110100111;
		16'b0111010011100010: color_data = 12'b001110100111;
		16'b0111010011110110: color_data = 12'b001110100111;
		16'b0111010011110111: color_data = 12'b001110100111;
		16'b0111010011111000: color_data = 12'b001110100111;
		16'b0111010011111001: color_data = 12'b001110100111;
		16'b0111010011111010: color_data = 12'b001110100111;
		16'b0111010011111011: color_data = 12'b001110100111;
		16'b0111010011111100: color_data = 12'b001110100111;
		16'b0111010011111101: color_data = 12'b001110100111;
		16'b0111010011111110: color_data = 12'b001110100111;
		16'b0111010011111111: color_data = 12'b001110100111;
		16'b0111010100000000: color_data = 12'b001110100111;
		16'b0111010100000001: color_data = 12'b001110100111;
		16'b0111010100011010: color_data = 12'b001110100111;
		16'b0111010100011011: color_data = 12'b001110100111;
		16'b0111010100011100: color_data = 12'b001110100111;
		16'b0111010100011101: color_data = 12'b001110100111;
		16'b0111010100011110: color_data = 12'b001110100111;
		16'b0111010100011111: color_data = 12'b001110100111;
		16'b0111010100100000: color_data = 12'b001110100111;
		16'b0111010100100001: color_data = 12'b001110100111;
		16'b0111010100100010: color_data = 12'b001110100111;
		16'b0111010100100011: color_data = 12'b001110100111;
		16'b0111010100100100: color_data = 12'b001110100111;
		16'b0111010100100101: color_data = 12'b001110100111;
		16'b0111010100100110: color_data = 12'b001110100111;
		16'b0111010100101101: color_data = 12'b001110100111;
		16'b0111010100101110: color_data = 12'b001110100111;
		16'b0111010100101111: color_data = 12'b001110100111;
		16'b0111010100110000: color_data = 12'b001110100111;
		16'b0111010100110001: color_data = 12'b001110100111;
		16'b0111010100110010: color_data = 12'b001110100111;
		16'b0111010100110011: color_data = 12'b001110100111;
		16'b0111010100110100: color_data = 12'b001110100111;
		16'b0111010100110101: color_data = 12'b001110100111;
		16'b0111010100110110: color_data = 12'b001110100111;
		16'b0111010100110111: color_data = 12'b001110100111;
		16'b0111010100111000: color_data = 12'b001110100111;
		16'b0111010101000101: color_data = 12'b001110100111;
		16'b0111010101000110: color_data = 12'b001110100111;
		16'b0111010101000111: color_data = 12'b001110100111;
		16'b0111010101001000: color_data = 12'b001110100111;
		16'b0111010101001001: color_data = 12'b001110100111;
		16'b0111010101001010: color_data = 12'b001110100111;
		16'b0111010101001011: color_data = 12'b001110100111;
		16'b0111010101001100: color_data = 12'b001110100111;
		16'b0111010101001101: color_data = 12'b001110100111;
		16'b0111010101001110: color_data = 12'b001110100111;
		16'b0111010101001111: color_data = 12'b001110100111;
		16'b0111010101010000: color_data = 12'b001110100111;
		16'b0111010101010001: color_data = 12'b001110100111;
		16'b0111010101011000: color_data = 12'b001110100111;
		16'b0111010101011001: color_data = 12'b001110100111;
		16'b0111010101011010: color_data = 12'b001110100111;
		16'b0111010101011011: color_data = 12'b001110100111;
		16'b0111010101011100: color_data = 12'b001110100111;
		16'b0111010101011101: color_data = 12'b001110100111;
		16'b0111010101011110: color_data = 12'b001110100111;
		16'b0111010101011111: color_data = 12'b001110100111;
		16'b0111010101100000: color_data = 12'b001110100111;
		16'b0111010101100001: color_data = 12'b001110100111;
		16'b0111010101100010: color_data = 12'b001110100111;
		16'b0111010101100011: color_data = 12'b001110100111;
		16'b0111010101110000: color_data = 12'b001110100111;
		16'b0111010101110001: color_data = 12'b001110100111;
		16'b0111010101110010: color_data = 12'b001110100111;
		16'b0111010101110011: color_data = 12'b001110100111;
		16'b0111010101110100: color_data = 12'b001110100111;
		16'b0111010101110101: color_data = 12'b001110100111;
		16'b0111010101110110: color_data = 12'b001110100111;
		16'b0111010101110111: color_data = 12'b001110100111;
		16'b0111010101111000: color_data = 12'b001110100111;
		16'b0111010101111001: color_data = 12'b001110100111;
		16'b0111010101111010: color_data = 12'b001110100111;
		16'b0111010101111011: color_data = 12'b001110100111;
		16'b0111011000000000: color_data = 12'b001110100111;
		16'b0111011000000001: color_data = 12'b001110100111;
		16'b0111011000000010: color_data = 12'b001110100111;
		16'b0111011000000011: color_data = 12'b001110100111;
		16'b0111011000000100: color_data = 12'b001110100111;
		16'b0111011000000101: color_data = 12'b001110100111;
		16'b0111011000000110: color_data = 12'b001110100111;
		16'b0111011000000111: color_data = 12'b001110100111;
		16'b0111011000001000: color_data = 12'b001110100111;
		16'b0111011000001001: color_data = 12'b001110100111;
		16'b0111011000001010: color_data = 12'b001110100111;
		16'b0111011000001011: color_data = 12'b001110100111;
		16'b0111011000001100: color_data = 12'b001110100111;
		16'b0111011000101011: color_data = 12'b001110100111;
		16'b0111011000101100: color_data = 12'b001110100111;
		16'b0111011000101101: color_data = 12'b001110100111;
		16'b0111011000101110: color_data = 12'b001110100111;
		16'b0111011000101111: color_data = 12'b001110100111;
		16'b0111011000110000: color_data = 12'b001110100111;
		16'b0111011000110001: color_data = 12'b001110100111;
		16'b0111011000110010: color_data = 12'b001110100111;
		16'b0111011000110011: color_data = 12'b001110100111;
		16'b0111011000110100: color_data = 12'b001110100111;
		16'b0111011000110101: color_data = 12'b001110100111;
		16'b0111011000110110: color_data = 12'b001110100111;
		16'b0111011000110111: color_data = 12'b001110100111;
		16'b0111011000111000: color_data = 12'b001110100111;
		16'b0111011000111001: color_data = 12'b001110100111;
		16'b0111011000111010: color_data = 12'b001110100111;
		16'b0111011000111011: color_data = 12'b001110100111;
		16'b0111011000111100: color_data = 12'b001110100111;
		16'b0111011000111101: color_data = 12'b001110100111;
		16'b0111011000111110: color_data = 12'b001110100111;
		16'b0111011000111111: color_data = 12'b001110100111;
		16'b0111011001000000: color_data = 12'b001110100111;
		16'b0111011001000001: color_data = 12'b001110100111;
		16'b0111011001000010: color_data = 12'b001110100111;
		16'b0111011001000011: color_data = 12'b001110100111;
		16'b0111011001000100: color_data = 12'b001110100111;
		16'b0111011001000101: color_data = 12'b001110100111;
		16'b0111011001000110: color_data = 12'b001110100111;
		16'b0111011001000111: color_data = 12'b001110100111;
		16'b0111011001001000: color_data = 12'b001110100111;
		16'b0111011001001001: color_data = 12'b001110100111;
		16'b0111011001001010: color_data = 12'b001110100111;
		16'b0111011001001011: color_data = 12'b001110100111;
		16'b0111011001001100: color_data = 12'b001110100111;
		16'b0111011001001101: color_data = 12'b001110100111;
		16'b0111011001001110: color_data = 12'b001110100111;
		16'b0111011001001111: color_data = 12'b001110100111;
		16'b0111011001011100: color_data = 12'b001110100111;
		16'b0111011001011101: color_data = 12'b001110100111;
		16'b0111011001011110: color_data = 12'b001110100111;
		16'b0111011001011111: color_data = 12'b001110100111;
		16'b0111011001100000: color_data = 12'b001110100111;
		16'b0111011001100001: color_data = 12'b001110100111;
		16'b0111011001100010: color_data = 12'b001110100111;
		16'b0111011001100011: color_data = 12'b001110100111;
		16'b0111011001100100: color_data = 12'b001110100111;
		16'b0111011001100101: color_data = 12'b001110100111;
		16'b0111011001100110: color_data = 12'b001110100111;
		16'b0111011001100111: color_data = 12'b001110100111;
		16'b0111011001101000: color_data = 12'b001110100111;
		16'b0111011001110101: color_data = 12'b001110100111;
		16'b0111011001110110: color_data = 12'b001110100111;
		16'b0111011001110111: color_data = 12'b001110100111;
		16'b0111011001111000: color_data = 12'b001110100111;
		16'b0111011001111001: color_data = 12'b001110100111;
		16'b0111011001111010: color_data = 12'b001110100111;
		16'b0111011001111011: color_data = 12'b001110100111;
		16'b0111011001111100: color_data = 12'b001110100111;
		16'b0111011001111101: color_data = 12'b001110100111;
		16'b0111011001111110: color_data = 12'b001110100111;
		16'b0111011001111111: color_data = 12'b001110100111;
		16'b0111011010000000: color_data = 12'b001110100111;
		16'b0111011010001101: color_data = 12'b001110100111;
		16'b0111011010001110: color_data = 12'b001110100111;
		16'b0111011010001111: color_data = 12'b001110100111;
		16'b0111011010010000: color_data = 12'b001110100111;
		16'b0111011010010001: color_data = 12'b001110100111;
		16'b0111011010010010: color_data = 12'b001110100111;
		16'b0111011010010011: color_data = 12'b001110100111;
		16'b0111011010010100: color_data = 12'b001110100111;
		16'b0111011010010101: color_data = 12'b001110100111;
		16'b0111011010010110: color_data = 12'b001110100111;
		16'b0111011010010111: color_data = 12'b001110100111;
		16'b0111011010011000: color_data = 12'b001110100111;
		16'b0111011010011001: color_data = 12'b001110100111;
		16'b0111011010100000: color_data = 12'b001110100111;
		16'b0111011010100001: color_data = 12'b001110100111;
		16'b0111011010100010: color_data = 12'b001110100111;
		16'b0111011010100011: color_data = 12'b001110100111;
		16'b0111011010100100: color_data = 12'b001110100111;
		16'b0111011010100101: color_data = 12'b001110100111;
		16'b0111011010100110: color_data = 12'b001110100111;
		16'b0111011010100111: color_data = 12'b001110100111;
		16'b0111011010101000: color_data = 12'b001110100111;
		16'b0111011010101001: color_data = 12'b001110100111;
		16'b0111011010101010: color_data = 12'b001110100111;
		16'b0111011010101011: color_data = 12'b001110100111;
		16'b0111011010111000: color_data = 12'b001110100111;
		16'b0111011010111001: color_data = 12'b001110100111;
		16'b0111011010111010: color_data = 12'b001110100111;
		16'b0111011010111011: color_data = 12'b001110100111;
		16'b0111011010111100: color_data = 12'b001110100111;
		16'b0111011010111101: color_data = 12'b001110100111;
		16'b0111011010111110: color_data = 12'b001110100111;
		16'b0111011010111111: color_data = 12'b001110100111;
		16'b0111011011000000: color_data = 12'b001110100111;
		16'b0111011011000001: color_data = 12'b001110100111;
		16'b0111011011000010: color_data = 12'b001110100111;
		16'b0111011011000011: color_data = 12'b001110100111;
		16'b0111011011000100: color_data = 12'b001110100111;
		16'b0111011011001011: color_data = 12'b001110100111;
		16'b0111011011001100: color_data = 12'b001110100111;
		16'b0111011011001101: color_data = 12'b001110100111;
		16'b0111011011001110: color_data = 12'b001110100111;
		16'b0111011011001111: color_data = 12'b001110100111;
		16'b0111011011010000: color_data = 12'b001110100111;
		16'b0111011011010001: color_data = 12'b001110100111;
		16'b0111011011010010: color_data = 12'b001110100111;
		16'b0111011011010011: color_data = 12'b001110100111;
		16'b0111011011010100: color_data = 12'b001110100111;
		16'b0111011011010101: color_data = 12'b001110100111;
		16'b0111011011010110: color_data = 12'b001110100111;
		16'b0111011011010111: color_data = 12'b001110100111;
		16'b0111011011011000: color_data = 12'b001110100111;
		16'b0111011011011001: color_data = 12'b001110100111;
		16'b0111011011011010: color_data = 12'b001110100111;
		16'b0111011011011011: color_data = 12'b001110100111;
		16'b0111011011011100: color_data = 12'b001110100111;
		16'b0111011011011101: color_data = 12'b001110100111;
		16'b0111011011011110: color_data = 12'b001110100111;
		16'b0111011011011111: color_data = 12'b001110100111;
		16'b0111011011100000: color_data = 12'b001110100111;
		16'b0111011011100001: color_data = 12'b001110100111;
		16'b0111011011100010: color_data = 12'b001110100111;
		16'b0111011011110110: color_data = 12'b001110100111;
		16'b0111011011110111: color_data = 12'b001110100111;
		16'b0111011011111000: color_data = 12'b001110100111;
		16'b0111011011111001: color_data = 12'b001110100111;
		16'b0111011011111010: color_data = 12'b001110100111;
		16'b0111011011111011: color_data = 12'b001110100111;
		16'b0111011011111100: color_data = 12'b001110100111;
		16'b0111011011111101: color_data = 12'b001110100111;
		16'b0111011011111110: color_data = 12'b001110100111;
		16'b0111011011111111: color_data = 12'b001110100111;
		16'b0111011100000000: color_data = 12'b001110100111;
		16'b0111011100000001: color_data = 12'b001110100111;
		16'b0111011100011010: color_data = 12'b001110100111;
		16'b0111011100011011: color_data = 12'b001110100111;
		16'b0111011100011100: color_data = 12'b001110100111;
		16'b0111011100011101: color_data = 12'b001110100111;
		16'b0111011100011110: color_data = 12'b001110100111;
		16'b0111011100011111: color_data = 12'b001110100111;
		16'b0111011100100000: color_data = 12'b001110100111;
		16'b0111011100100001: color_data = 12'b001110100111;
		16'b0111011100100010: color_data = 12'b001110100111;
		16'b0111011100100011: color_data = 12'b001110100111;
		16'b0111011100100100: color_data = 12'b001110100111;
		16'b0111011100100101: color_data = 12'b001110100111;
		16'b0111011100100110: color_data = 12'b001110100111;
		16'b0111011100101101: color_data = 12'b001110100111;
		16'b0111011100101110: color_data = 12'b001110100111;
		16'b0111011100101111: color_data = 12'b001110100111;
		16'b0111011100110000: color_data = 12'b001110100111;
		16'b0111011100110001: color_data = 12'b001110100111;
		16'b0111011100110010: color_data = 12'b001110100111;
		16'b0111011100110011: color_data = 12'b001110100111;
		16'b0111011100110100: color_data = 12'b001110100111;
		16'b0111011100110101: color_data = 12'b001110100111;
		16'b0111011100110110: color_data = 12'b001110100111;
		16'b0111011100110111: color_data = 12'b001110100111;
		16'b0111011100111000: color_data = 12'b001110100111;
		16'b0111011101000101: color_data = 12'b001110100111;
		16'b0111011101000110: color_data = 12'b001110100111;
		16'b0111011101000111: color_data = 12'b001110100111;
		16'b0111011101001000: color_data = 12'b001110100111;
		16'b0111011101001001: color_data = 12'b001110100111;
		16'b0111011101001010: color_data = 12'b001110100111;
		16'b0111011101001011: color_data = 12'b001110100111;
		16'b0111011101001100: color_data = 12'b001110100111;
		16'b0111011101001101: color_data = 12'b001110100111;
		16'b0111011101001110: color_data = 12'b001110100111;
		16'b0111011101001111: color_data = 12'b001110100111;
		16'b0111011101010000: color_data = 12'b001110100111;
		16'b0111011101010001: color_data = 12'b001110100111;
		16'b0111011101011000: color_data = 12'b001110100111;
		16'b0111011101011001: color_data = 12'b001110100111;
		16'b0111011101011010: color_data = 12'b001110100111;
		16'b0111011101011011: color_data = 12'b001110100111;
		16'b0111011101011100: color_data = 12'b001110100111;
		16'b0111011101011101: color_data = 12'b001110100111;
		16'b0111011101011110: color_data = 12'b001110100111;
		16'b0111011101011111: color_data = 12'b001110100111;
		16'b0111011101100000: color_data = 12'b001110100111;
		16'b0111011101100001: color_data = 12'b001110100111;
		16'b0111011101100010: color_data = 12'b001110100111;
		16'b0111011101100011: color_data = 12'b001110100111;
		16'b0111011101110000: color_data = 12'b001110100111;
		16'b0111011101110001: color_data = 12'b001110100111;
		16'b0111011101110010: color_data = 12'b001110100111;
		16'b0111011101110011: color_data = 12'b001110100111;
		16'b0111011101110100: color_data = 12'b001110100111;
		16'b0111011101110101: color_data = 12'b001110100111;
		16'b0111011101110110: color_data = 12'b001110100111;
		16'b0111011101110111: color_data = 12'b001110100111;
		16'b0111011101111000: color_data = 12'b001110100111;
		16'b0111011101111001: color_data = 12'b001110100111;
		16'b0111011101111010: color_data = 12'b001110100111;
		16'b0111011101111011: color_data = 12'b001110100111;
		16'b0111100000000000: color_data = 12'b001110100111;
		16'b0111100000000001: color_data = 12'b001110100111;
		16'b0111100000000010: color_data = 12'b001110100111;
		16'b0111100000000011: color_data = 12'b001110100111;
		16'b0111100000000100: color_data = 12'b001110100111;
		16'b0111100000000101: color_data = 12'b001110100111;
		16'b0111100000000110: color_data = 12'b001110100111;
		16'b0111100000000111: color_data = 12'b001110100111;
		16'b0111100000001000: color_data = 12'b001110100111;
		16'b0111100000001001: color_data = 12'b001110100111;
		16'b0111100000001010: color_data = 12'b001110100111;
		16'b0111100000001011: color_data = 12'b001110100111;
		16'b0111100000001100: color_data = 12'b001110100111;
		16'b0111100000101011: color_data = 12'b001110100111;
		16'b0111100000101100: color_data = 12'b001110100111;
		16'b0111100000101101: color_data = 12'b001110100111;
		16'b0111100000101110: color_data = 12'b001110100111;
		16'b0111100000101111: color_data = 12'b001110100111;
		16'b0111100000110000: color_data = 12'b001110100111;
		16'b0111100000110001: color_data = 12'b001110100111;
		16'b0111100000110010: color_data = 12'b001110100111;
		16'b0111100000110011: color_data = 12'b001110100111;
		16'b0111100000110100: color_data = 12'b001110100111;
		16'b0111100000110101: color_data = 12'b001110100111;
		16'b0111100000110110: color_data = 12'b001110100111;
		16'b0111100000110111: color_data = 12'b001110100111;
		16'b0111100000111000: color_data = 12'b001110100111;
		16'b0111100000111001: color_data = 12'b001110100111;
		16'b0111100000111010: color_data = 12'b001110100111;
		16'b0111100000111011: color_data = 12'b001110100111;
		16'b0111100000111100: color_data = 12'b001110100111;
		16'b0111100000111101: color_data = 12'b001110100111;
		16'b0111100000111110: color_data = 12'b001110100111;
		16'b0111100000111111: color_data = 12'b001110100111;
		16'b0111100001000000: color_data = 12'b001110100111;
		16'b0111100001000001: color_data = 12'b001110100111;
		16'b0111100001000010: color_data = 12'b001110100111;
		16'b0111100001000011: color_data = 12'b001110100111;
		16'b0111100001000100: color_data = 12'b001110100111;
		16'b0111100001000101: color_data = 12'b001110100111;
		16'b0111100001000110: color_data = 12'b001110100111;
		16'b0111100001000111: color_data = 12'b001110100111;
		16'b0111100001001000: color_data = 12'b001110100111;
		16'b0111100001001001: color_data = 12'b001110100111;
		16'b0111100001001010: color_data = 12'b001110100111;
		16'b0111100001001011: color_data = 12'b001110100111;
		16'b0111100001001100: color_data = 12'b001110100111;
		16'b0111100001001101: color_data = 12'b001110100111;
		16'b0111100001001110: color_data = 12'b001110100111;
		16'b0111100001001111: color_data = 12'b001110100111;
		16'b0111100001011100: color_data = 12'b001110100111;
		16'b0111100001011101: color_data = 12'b001110100111;
		16'b0111100001011110: color_data = 12'b001110100111;
		16'b0111100001011111: color_data = 12'b001110100111;
		16'b0111100001100000: color_data = 12'b001110100111;
		16'b0111100001100001: color_data = 12'b001110100111;
		16'b0111100001100010: color_data = 12'b001110100111;
		16'b0111100001100011: color_data = 12'b001110100111;
		16'b0111100001100100: color_data = 12'b001110100111;
		16'b0111100001100101: color_data = 12'b001110100111;
		16'b0111100001100110: color_data = 12'b001110100111;
		16'b0111100001100111: color_data = 12'b001110100111;
		16'b0111100001101000: color_data = 12'b001110100111;
		16'b0111100001110101: color_data = 12'b001110100111;
		16'b0111100001110110: color_data = 12'b001110100111;
		16'b0111100001110111: color_data = 12'b001110100111;
		16'b0111100001111000: color_data = 12'b001110100111;
		16'b0111100001111001: color_data = 12'b001110100111;
		16'b0111100001111010: color_data = 12'b001110100111;
		16'b0111100001111011: color_data = 12'b001110100111;
		16'b0111100001111100: color_data = 12'b001110100111;
		16'b0111100001111101: color_data = 12'b001110100111;
		16'b0111100001111110: color_data = 12'b001110100111;
		16'b0111100001111111: color_data = 12'b001110100111;
		16'b0111100010000000: color_data = 12'b001110100111;
		16'b0111100010001101: color_data = 12'b001110100111;
		16'b0111100010001110: color_data = 12'b001110100111;
		16'b0111100010001111: color_data = 12'b001110100111;
		16'b0111100010010000: color_data = 12'b001110100111;
		16'b0111100010010001: color_data = 12'b001110100111;
		16'b0111100010010010: color_data = 12'b001110100111;
		16'b0111100010010011: color_data = 12'b001110100111;
		16'b0111100010010100: color_data = 12'b001110100111;
		16'b0111100010010101: color_data = 12'b001110100111;
		16'b0111100010010110: color_data = 12'b001110100111;
		16'b0111100010010111: color_data = 12'b001110100111;
		16'b0111100010011000: color_data = 12'b001110100111;
		16'b0111100010011001: color_data = 12'b001110100111;
		16'b0111100010100000: color_data = 12'b001110100111;
		16'b0111100010100001: color_data = 12'b001110100111;
		16'b0111100010100010: color_data = 12'b001110100111;
		16'b0111100010100011: color_data = 12'b001110100111;
		16'b0111100010100100: color_data = 12'b001110100111;
		16'b0111100010100101: color_data = 12'b001110100111;
		16'b0111100010100110: color_data = 12'b001110100111;
		16'b0111100010100111: color_data = 12'b001110100111;
		16'b0111100010101000: color_data = 12'b001110100111;
		16'b0111100010101001: color_data = 12'b001110100111;
		16'b0111100010101010: color_data = 12'b001110100111;
		16'b0111100010101011: color_data = 12'b001110100111;
		16'b0111100010111000: color_data = 12'b001110100111;
		16'b0111100010111001: color_data = 12'b001110100111;
		16'b0111100010111010: color_data = 12'b001110100111;
		16'b0111100010111011: color_data = 12'b001110100111;
		16'b0111100010111100: color_data = 12'b001110100111;
		16'b0111100010111101: color_data = 12'b001110100111;
		16'b0111100010111110: color_data = 12'b001110100111;
		16'b0111100010111111: color_data = 12'b001110100111;
		16'b0111100011000000: color_data = 12'b001110100111;
		16'b0111100011000001: color_data = 12'b001110100111;
		16'b0111100011000010: color_data = 12'b001110100111;
		16'b0111100011000011: color_data = 12'b001110100111;
		16'b0111100011000100: color_data = 12'b001110100111;
		16'b0111100011001011: color_data = 12'b001110100111;
		16'b0111100011001100: color_data = 12'b001110100111;
		16'b0111100011001101: color_data = 12'b001110100111;
		16'b0111100011001110: color_data = 12'b001110100111;
		16'b0111100011001111: color_data = 12'b001110100111;
		16'b0111100011010000: color_data = 12'b001110100111;
		16'b0111100011010001: color_data = 12'b001110100111;
		16'b0111100011010010: color_data = 12'b001110100111;
		16'b0111100011010011: color_data = 12'b001110100111;
		16'b0111100011010100: color_data = 12'b001110100111;
		16'b0111100011010101: color_data = 12'b001110100111;
		16'b0111100011010110: color_data = 12'b001110100111;
		16'b0111100011010111: color_data = 12'b001110100111;
		16'b0111100011011000: color_data = 12'b001110100111;
		16'b0111100011011001: color_data = 12'b001110100111;
		16'b0111100011011010: color_data = 12'b001110100111;
		16'b0111100011011011: color_data = 12'b001110100111;
		16'b0111100011011100: color_data = 12'b001110100111;
		16'b0111100011011101: color_data = 12'b001110100111;
		16'b0111100011011110: color_data = 12'b001110100111;
		16'b0111100011011111: color_data = 12'b001110100111;
		16'b0111100011100000: color_data = 12'b001110100111;
		16'b0111100011100001: color_data = 12'b001110100111;
		16'b0111100011100010: color_data = 12'b001110100111;
		16'b0111100011110110: color_data = 12'b001110100111;
		16'b0111100011110111: color_data = 12'b001110100111;
		16'b0111100011111000: color_data = 12'b001110100111;
		16'b0111100011111001: color_data = 12'b001110100111;
		16'b0111100011111010: color_data = 12'b001110100111;
		16'b0111100011111011: color_data = 12'b001110100111;
		16'b0111100011111100: color_data = 12'b001110100111;
		16'b0111100011111101: color_data = 12'b001110100111;
		16'b0111100011111110: color_data = 12'b001110100111;
		16'b0111100011111111: color_data = 12'b001110100111;
		16'b0111100100000000: color_data = 12'b001110100111;
		16'b0111100100000001: color_data = 12'b001110100111;
		16'b0111100100011010: color_data = 12'b001110100111;
		16'b0111100100011011: color_data = 12'b001110100111;
		16'b0111100100011100: color_data = 12'b001110100111;
		16'b0111100100011101: color_data = 12'b001110100111;
		16'b0111100100011110: color_data = 12'b001110100111;
		16'b0111100100011111: color_data = 12'b001110100111;
		16'b0111100100100000: color_data = 12'b001110100111;
		16'b0111100100100001: color_data = 12'b001110100111;
		16'b0111100100100010: color_data = 12'b001110100111;
		16'b0111100100100011: color_data = 12'b001110100111;
		16'b0111100100100100: color_data = 12'b001110100111;
		16'b0111100100100101: color_data = 12'b001110100111;
		16'b0111100100100110: color_data = 12'b001110100111;
		16'b0111100100101101: color_data = 12'b001110100111;
		16'b0111100100101110: color_data = 12'b001110100111;
		16'b0111100100101111: color_data = 12'b001110100111;
		16'b0111100100110000: color_data = 12'b001110100111;
		16'b0111100100110001: color_data = 12'b001110100111;
		16'b0111100100110010: color_data = 12'b001110100111;
		16'b0111100100110011: color_data = 12'b001110100111;
		16'b0111100100110100: color_data = 12'b001110100111;
		16'b0111100100110101: color_data = 12'b001110100111;
		16'b0111100100110110: color_data = 12'b001110100111;
		16'b0111100100110111: color_data = 12'b001110100111;
		16'b0111100100111000: color_data = 12'b001110100111;
		16'b0111100101000101: color_data = 12'b001110100111;
		16'b0111100101000110: color_data = 12'b001110100111;
		16'b0111100101000111: color_data = 12'b001110100111;
		16'b0111100101001000: color_data = 12'b001110100111;
		16'b0111100101001001: color_data = 12'b001110100111;
		16'b0111100101001010: color_data = 12'b001110100111;
		16'b0111100101001011: color_data = 12'b001110100111;
		16'b0111100101001100: color_data = 12'b001110100111;
		16'b0111100101001101: color_data = 12'b001110100111;
		16'b0111100101001110: color_data = 12'b001110100111;
		16'b0111100101001111: color_data = 12'b001110100111;
		16'b0111100101010000: color_data = 12'b001110100111;
		16'b0111100101010001: color_data = 12'b001110100111;
		16'b0111100101011000: color_data = 12'b001110100111;
		16'b0111100101011001: color_data = 12'b001110100111;
		16'b0111100101011010: color_data = 12'b001110100111;
		16'b0111100101011011: color_data = 12'b001110100111;
		16'b0111100101011100: color_data = 12'b001110100111;
		16'b0111100101011101: color_data = 12'b001110100111;
		16'b0111100101011110: color_data = 12'b001110100111;
		16'b0111100101011111: color_data = 12'b001110100111;
		16'b0111100101100000: color_data = 12'b001110100111;
		16'b0111100101100001: color_data = 12'b001110100111;
		16'b0111100101100010: color_data = 12'b001110100111;
		16'b0111100101100011: color_data = 12'b001110100111;
		16'b0111100101110000: color_data = 12'b001110100111;
		16'b0111100101110001: color_data = 12'b001110100111;
		16'b0111100101110010: color_data = 12'b001110100111;
		16'b0111100101110011: color_data = 12'b001110100111;
		16'b0111100101110100: color_data = 12'b001110100111;
		16'b0111100101110101: color_data = 12'b001110100111;
		16'b0111100101110110: color_data = 12'b001110100111;
		16'b0111100101110111: color_data = 12'b001110100111;
		16'b0111100101111000: color_data = 12'b001110100111;
		16'b0111100101111001: color_data = 12'b001110100111;
		16'b0111100101111010: color_data = 12'b001110100111;
		16'b0111100101111011: color_data = 12'b001110100111;
		16'b0111101000000000: color_data = 12'b001110100111;
		16'b0111101000000001: color_data = 12'b001110100111;
		16'b0111101000000010: color_data = 12'b001110100111;
		16'b0111101000000011: color_data = 12'b001110100111;
		16'b0111101000000100: color_data = 12'b001110100111;
		16'b0111101000000101: color_data = 12'b001110100111;
		16'b0111101000000110: color_data = 12'b001110100111;
		16'b0111101000000111: color_data = 12'b001110100111;
		16'b0111101000001000: color_data = 12'b001110100111;
		16'b0111101000001001: color_data = 12'b001110100111;
		16'b0111101000001010: color_data = 12'b001110100111;
		16'b0111101000001011: color_data = 12'b001110100111;
		16'b0111101000001100: color_data = 12'b001110100111;
		16'b0111101000101011: color_data = 12'b001110100111;
		16'b0111101000101100: color_data = 12'b001110100111;
		16'b0111101000101101: color_data = 12'b001110100111;
		16'b0111101000101110: color_data = 12'b001110100111;
		16'b0111101000101111: color_data = 12'b001110100111;
		16'b0111101000110000: color_data = 12'b001110100111;
		16'b0111101000110001: color_data = 12'b001110100111;
		16'b0111101000110010: color_data = 12'b001110100111;
		16'b0111101000110011: color_data = 12'b001110100111;
		16'b0111101000110100: color_data = 12'b001110100111;
		16'b0111101000110101: color_data = 12'b001110100111;
		16'b0111101000110110: color_data = 12'b001110100111;
		16'b0111101000110111: color_data = 12'b001110100111;
		16'b0111101000111000: color_data = 12'b001110100111;
		16'b0111101000111001: color_data = 12'b001110100111;
		16'b0111101000111010: color_data = 12'b001110100111;
		16'b0111101000111011: color_data = 12'b001110100111;
		16'b0111101000111100: color_data = 12'b001110100111;
		16'b0111101000111101: color_data = 12'b001110100111;
		16'b0111101000111110: color_data = 12'b001110100111;
		16'b0111101000111111: color_data = 12'b001110100111;
		16'b0111101001000000: color_data = 12'b001110100111;
		16'b0111101001000001: color_data = 12'b001110100111;
		16'b0111101001000010: color_data = 12'b001110100111;
		16'b0111101001000011: color_data = 12'b001110100111;
		16'b0111101001000100: color_data = 12'b001110100111;
		16'b0111101001000101: color_data = 12'b001110100111;
		16'b0111101001000110: color_data = 12'b001110100111;
		16'b0111101001000111: color_data = 12'b001110100111;
		16'b0111101001001000: color_data = 12'b001110100111;
		16'b0111101001001001: color_data = 12'b001110100111;
		16'b0111101001001010: color_data = 12'b001110100111;
		16'b0111101001001011: color_data = 12'b001110100111;
		16'b0111101001001100: color_data = 12'b001110100111;
		16'b0111101001001101: color_data = 12'b001110100111;
		16'b0111101001001110: color_data = 12'b001110100111;
		16'b0111101001001111: color_data = 12'b001110100111;
		16'b0111101001011100: color_data = 12'b001110100111;
		16'b0111101001011101: color_data = 12'b001110100111;
		16'b0111101001011110: color_data = 12'b001110100111;
		16'b0111101001011111: color_data = 12'b001110100111;
		16'b0111101001100000: color_data = 12'b001110100111;
		16'b0111101001100001: color_data = 12'b001110100111;
		16'b0111101001100010: color_data = 12'b001110100111;
		16'b0111101001100011: color_data = 12'b001110100111;
		16'b0111101001100100: color_data = 12'b001110100111;
		16'b0111101001100101: color_data = 12'b001110100111;
		16'b0111101001100110: color_data = 12'b001110100111;
		16'b0111101001100111: color_data = 12'b001110100111;
		16'b0111101001101000: color_data = 12'b001110100111;
		16'b0111101001110101: color_data = 12'b001110100111;
		16'b0111101001110110: color_data = 12'b001110100111;
		16'b0111101001110111: color_data = 12'b001110100111;
		16'b0111101001111000: color_data = 12'b001110100111;
		16'b0111101001111001: color_data = 12'b001110100111;
		16'b0111101001111010: color_data = 12'b001110100111;
		16'b0111101001111011: color_data = 12'b001110100111;
		16'b0111101001111100: color_data = 12'b001110100111;
		16'b0111101001111101: color_data = 12'b001110100111;
		16'b0111101001111110: color_data = 12'b001110100111;
		16'b0111101001111111: color_data = 12'b001110100111;
		16'b0111101010000000: color_data = 12'b001110100111;
		16'b0111101010001101: color_data = 12'b001110100111;
		16'b0111101010001110: color_data = 12'b001110100111;
		16'b0111101010001111: color_data = 12'b001110100111;
		16'b0111101010010000: color_data = 12'b001110100111;
		16'b0111101010010001: color_data = 12'b001110100111;
		16'b0111101010010010: color_data = 12'b001110100111;
		16'b0111101010010011: color_data = 12'b001110100111;
		16'b0111101010010100: color_data = 12'b001110100111;
		16'b0111101010010101: color_data = 12'b001110100111;
		16'b0111101010010110: color_data = 12'b001110100111;
		16'b0111101010010111: color_data = 12'b001110100111;
		16'b0111101010011000: color_data = 12'b001110100111;
		16'b0111101010011001: color_data = 12'b001110100111;
		16'b0111101010100000: color_data = 12'b001110100111;
		16'b0111101010100001: color_data = 12'b001110100111;
		16'b0111101010100010: color_data = 12'b001110100111;
		16'b0111101010100011: color_data = 12'b001110100111;
		16'b0111101010100100: color_data = 12'b001110100111;
		16'b0111101010100101: color_data = 12'b001110100111;
		16'b0111101010100110: color_data = 12'b001110100111;
		16'b0111101010100111: color_data = 12'b001110100111;
		16'b0111101010101000: color_data = 12'b001110100111;
		16'b0111101010101001: color_data = 12'b001110100111;
		16'b0111101010101010: color_data = 12'b001110100111;
		16'b0111101010101011: color_data = 12'b001110100111;
		16'b0111101010111000: color_data = 12'b001110100111;
		16'b0111101010111001: color_data = 12'b001110100111;
		16'b0111101010111010: color_data = 12'b001110100111;
		16'b0111101010111011: color_data = 12'b001110100111;
		16'b0111101010111100: color_data = 12'b001110100111;
		16'b0111101010111101: color_data = 12'b001110100111;
		16'b0111101010111110: color_data = 12'b001110100111;
		16'b0111101010111111: color_data = 12'b001110100111;
		16'b0111101011000000: color_data = 12'b001110100111;
		16'b0111101011000001: color_data = 12'b001110100111;
		16'b0111101011000010: color_data = 12'b001110100111;
		16'b0111101011000011: color_data = 12'b001110100111;
		16'b0111101011000100: color_data = 12'b001110100111;
		16'b0111101011001011: color_data = 12'b001110100111;
		16'b0111101011001100: color_data = 12'b001110100111;
		16'b0111101011001101: color_data = 12'b001110100111;
		16'b0111101011001110: color_data = 12'b001110100111;
		16'b0111101011001111: color_data = 12'b001110100111;
		16'b0111101011010000: color_data = 12'b001110100111;
		16'b0111101011010001: color_data = 12'b001110100111;
		16'b0111101011010010: color_data = 12'b001110100111;
		16'b0111101011010011: color_data = 12'b001110100111;
		16'b0111101011010100: color_data = 12'b001110100111;
		16'b0111101011010101: color_data = 12'b001110100111;
		16'b0111101011010110: color_data = 12'b001110100111;
		16'b0111101011010111: color_data = 12'b001110100111;
		16'b0111101011011000: color_data = 12'b001110100111;
		16'b0111101011011001: color_data = 12'b001110100111;
		16'b0111101011011010: color_data = 12'b001110100111;
		16'b0111101011011011: color_data = 12'b001110100111;
		16'b0111101011011100: color_data = 12'b001110100111;
		16'b0111101011011101: color_data = 12'b001110100111;
		16'b0111101011011110: color_data = 12'b001110100111;
		16'b0111101011011111: color_data = 12'b001110100111;
		16'b0111101011100000: color_data = 12'b001110100111;
		16'b0111101011100001: color_data = 12'b001110100111;
		16'b0111101011100010: color_data = 12'b001110100111;
		16'b0111101011110110: color_data = 12'b001110100111;
		16'b0111101011110111: color_data = 12'b001110100111;
		16'b0111101011111000: color_data = 12'b001110100111;
		16'b0111101011111001: color_data = 12'b001110100111;
		16'b0111101011111010: color_data = 12'b001110100111;
		16'b0111101011111011: color_data = 12'b001110100111;
		16'b0111101011111100: color_data = 12'b001110100111;
		16'b0111101011111101: color_data = 12'b001110100111;
		16'b0111101011111110: color_data = 12'b001110100111;
		16'b0111101011111111: color_data = 12'b001110100111;
		16'b0111101100000000: color_data = 12'b001110100111;
		16'b0111101100000001: color_data = 12'b001110100111;
		16'b0111101100011010: color_data = 12'b001110100111;
		16'b0111101100011011: color_data = 12'b001110100111;
		16'b0111101100011100: color_data = 12'b001110100111;
		16'b0111101100011101: color_data = 12'b001110100111;
		16'b0111101100011110: color_data = 12'b001110100111;
		16'b0111101100011111: color_data = 12'b001110100111;
		16'b0111101100100000: color_data = 12'b001110100111;
		16'b0111101100100001: color_data = 12'b001110100111;
		16'b0111101100100010: color_data = 12'b001110100111;
		16'b0111101100100011: color_data = 12'b001110100111;
		16'b0111101100100100: color_data = 12'b001110100111;
		16'b0111101100100101: color_data = 12'b001110100111;
		16'b0111101100100110: color_data = 12'b001110100111;
		16'b0111101100101101: color_data = 12'b001110100111;
		16'b0111101100101110: color_data = 12'b001110100111;
		16'b0111101100101111: color_data = 12'b001110100111;
		16'b0111101100110000: color_data = 12'b001110100111;
		16'b0111101100110001: color_data = 12'b001110100111;
		16'b0111101100110010: color_data = 12'b001110100111;
		16'b0111101100110011: color_data = 12'b001110100111;
		16'b0111101100110100: color_data = 12'b001110100111;
		16'b0111101100110101: color_data = 12'b001110100111;
		16'b0111101100110110: color_data = 12'b001110100111;
		16'b0111101100110111: color_data = 12'b001110100111;
		16'b0111101100111000: color_data = 12'b001110100111;
		16'b0111101101000101: color_data = 12'b001110100111;
		16'b0111101101000110: color_data = 12'b001110100111;
		16'b0111101101000111: color_data = 12'b001110100111;
		16'b0111101101001000: color_data = 12'b001110100111;
		16'b0111101101001001: color_data = 12'b001110100111;
		16'b0111101101001010: color_data = 12'b001110100111;
		16'b0111101101001011: color_data = 12'b001110100111;
		16'b0111101101001100: color_data = 12'b001110100111;
		16'b0111101101001101: color_data = 12'b001110100111;
		16'b0111101101001110: color_data = 12'b001110100111;
		16'b0111101101001111: color_data = 12'b001110100111;
		16'b0111101101010000: color_data = 12'b001110100111;
		16'b0111101101010001: color_data = 12'b001110100111;
		16'b0111101101011000: color_data = 12'b001110100111;
		16'b0111101101011001: color_data = 12'b001110100111;
		16'b0111101101011010: color_data = 12'b001110100111;
		16'b0111101101011011: color_data = 12'b001110100111;
		16'b0111101101011100: color_data = 12'b001110100111;
		16'b0111101101011101: color_data = 12'b001110100111;
		16'b0111101101011110: color_data = 12'b001110100111;
		16'b0111101101011111: color_data = 12'b001110100111;
		16'b0111101101100000: color_data = 12'b001110100111;
		16'b0111101101100001: color_data = 12'b001110100111;
		16'b0111101101100010: color_data = 12'b001110100111;
		16'b0111101101100011: color_data = 12'b001110100111;
		16'b0111101101110000: color_data = 12'b001110100111;
		16'b0111101101110001: color_data = 12'b001110100111;
		16'b0111101101110010: color_data = 12'b001110100111;
		16'b0111101101110011: color_data = 12'b001110100111;
		16'b0111101101110100: color_data = 12'b001110100111;
		16'b0111101101110101: color_data = 12'b001110100111;
		16'b0111101101110110: color_data = 12'b001110100111;
		16'b0111101101110111: color_data = 12'b001110100111;
		16'b0111101101111000: color_data = 12'b001110100111;
		16'b0111101101111001: color_data = 12'b001110100111;
		16'b0111101101111010: color_data = 12'b001110100111;
		16'b0111101101111011: color_data = 12'b001110100111;
		16'b0111110000000000: color_data = 12'b001110100111;
		16'b0111110000000001: color_data = 12'b001110100111;
		16'b0111110000000010: color_data = 12'b001110100111;
		16'b0111110000000011: color_data = 12'b001110100111;
		16'b0111110000000100: color_data = 12'b001110100111;
		16'b0111110000000101: color_data = 12'b001110100111;
		16'b0111110000000110: color_data = 12'b001110100111;
		16'b0111110000000111: color_data = 12'b001110100111;
		16'b0111110000001000: color_data = 12'b001110100111;
		16'b0111110000001001: color_data = 12'b001110100111;
		16'b0111110000001010: color_data = 12'b001110100111;
		16'b0111110000001011: color_data = 12'b001110100111;
		16'b0111110000001100: color_data = 12'b001110100111;
		16'b0111110000101011: color_data = 12'b001110100111;
		16'b0111110000101100: color_data = 12'b001110100111;
		16'b0111110000101101: color_data = 12'b001110100111;
		16'b0111110000101110: color_data = 12'b001110100111;
		16'b0111110000101111: color_data = 12'b001110100111;
		16'b0111110000110000: color_data = 12'b001110100111;
		16'b0111110000110001: color_data = 12'b001110100111;
		16'b0111110000110010: color_data = 12'b001110100111;
		16'b0111110000110011: color_data = 12'b001110100111;
		16'b0111110000110100: color_data = 12'b001110100111;
		16'b0111110000110101: color_data = 12'b001110100111;
		16'b0111110000110110: color_data = 12'b001110100111;
		16'b0111110000110111: color_data = 12'b001110100111;
		16'b0111110000111000: color_data = 12'b001110100111;
		16'b0111110000111001: color_data = 12'b001110100111;
		16'b0111110000111010: color_data = 12'b001110100111;
		16'b0111110000111011: color_data = 12'b001110100111;
		16'b0111110000111100: color_data = 12'b001110100111;
		16'b0111110000111101: color_data = 12'b001110100111;
		16'b0111110000111110: color_data = 12'b001110100111;
		16'b0111110000111111: color_data = 12'b001110100111;
		16'b0111110001000000: color_data = 12'b001110100111;
		16'b0111110001000001: color_data = 12'b001110100111;
		16'b0111110001000010: color_data = 12'b001110100111;
		16'b0111110001000011: color_data = 12'b001110100111;
		16'b0111110001000100: color_data = 12'b001110100111;
		16'b0111110001000101: color_data = 12'b001110100111;
		16'b0111110001000110: color_data = 12'b001110100111;
		16'b0111110001000111: color_data = 12'b001110100111;
		16'b0111110001001000: color_data = 12'b001110100111;
		16'b0111110001001001: color_data = 12'b001110100111;
		16'b0111110001001010: color_data = 12'b001110100111;
		16'b0111110001001011: color_data = 12'b001110100111;
		16'b0111110001001100: color_data = 12'b001110100111;
		16'b0111110001001101: color_data = 12'b001110100111;
		16'b0111110001001110: color_data = 12'b001110100111;
		16'b0111110001001111: color_data = 12'b001110100111;
		16'b0111110001011100: color_data = 12'b001110100111;
		16'b0111110001011101: color_data = 12'b001110100111;
		16'b0111110001011110: color_data = 12'b001110100111;
		16'b0111110001011111: color_data = 12'b001110100111;
		16'b0111110001100000: color_data = 12'b001110100111;
		16'b0111110001100001: color_data = 12'b001110100111;
		16'b0111110001100010: color_data = 12'b001110100111;
		16'b0111110001100011: color_data = 12'b001110100111;
		16'b0111110001100100: color_data = 12'b001110100111;
		16'b0111110001100101: color_data = 12'b001110100111;
		16'b0111110001100110: color_data = 12'b001110100111;
		16'b0111110001100111: color_data = 12'b001110100111;
		16'b0111110001101000: color_data = 12'b001110100111;
		16'b0111110001110101: color_data = 12'b001110100111;
		16'b0111110001110110: color_data = 12'b001110100111;
		16'b0111110001110111: color_data = 12'b001110100111;
		16'b0111110001111000: color_data = 12'b001110100111;
		16'b0111110001111001: color_data = 12'b001110100111;
		16'b0111110001111010: color_data = 12'b001110100111;
		16'b0111110001111011: color_data = 12'b001110100111;
		16'b0111110001111100: color_data = 12'b001110100111;
		16'b0111110001111101: color_data = 12'b001110100111;
		16'b0111110001111110: color_data = 12'b001110100111;
		16'b0111110001111111: color_data = 12'b001110100111;
		16'b0111110010000000: color_data = 12'b001110100111;
		16'b0111110010001101: color_data = 12'b001110100111;
		16'b0111110010001110: color_data = 12'b001110100111;
		16'b0111110010001111: color_data = 12'b001110100111;
		16'b0111110010010000: color_data = 12'b001110100111;
		16'b0111110010010001: color_data = 12'b001110100111;
		16'b0111110010010010: color_data = 12'b001110100111;
		16'b0111110010010011: color_data = 12'b001110100111;
		16'b0111110010010100: color_data = 12'b001110100111;
		16'b0111110010010101: color_data = 12'b001110100111;
		16'b0111110010010110: color_data = 12'b001110100111;
		16'b0111110010010111: color_data = 12'b001110100111;
		16'b0111110010011000: color_data = 12'b001110100111;
		16'b0111110010011001: color_data = 12'b001110100111;
		16'b0111110010100000: color_data = 12'b001110100111;
		16'b0111110010100001: color_data = 12'b001110100111;
		16'b0111110010100010: color_data = 12'b001110100111;
		16'b0111110010100011: color_data = 12'b001110100111;
		16'b0111110010100100: color_data = 12'b001110100111;
		16'b0111110010100101: color_data = 12'b001110100111;
		16'b0111110010100110: color_data = 12'b001110100111;
		16'b0111110010100111: color_data = 12'b001110100111;
		16'b0111110010101000: color_data = 12'b001110100111;
		16'b0111110010101001: color_data = 12'b001110100111;
		16'b0111110010101010: color_data = 12'b001110100111;
		16'b0111110010101011: color_data = 12'b001110100111;
		16'b0111110010111000: color_data = 12'b001110100111;
		16'b0111110010111001: color_data = 12'b001110100111;
		16'b0111110010111010: color_data = 12'b001110100111;
		16'b0111110010111011: color_data = 12'b001110100111;
		16'b0111110010111100: color_data = 12'b001110100111;
		16'b0111110010111101: color_data = 12'b001110100111;
		16'b0111110010111110: color_data = 12'b001110100111;
		16'b0111110010111111: color_data = 12'b001110100111;
		16'b0111110011000000: color_data = 12'b001110100111;
		16'b0111110011000001: color_data = 12'b001110100111;
		16'b0111110011000010: color_data = 12'b001110100111;
		16'b0111110011000011: color_data = 12'b001110100111;
		16'b0111110011000100: color_data = 12'b001110100111;
		16'b0111110011001011: color_data = 12'b001110100111;
		16'b0111110011001100: color_data = 12'b001110100111;
		16'b0111110011001101: color_data = 12'b001110100111;
		16'b0111110011001110: color_data = 12'b001110100111;
		16'b0111110011001111: color_data = 12'b001110100111;
		16'b0111110011010000: color_data = 12'b001110100111;
		16'b0111110011010001: color_data = 12'b001110100111;
		16'b0111110011010010: color_data = 12'b001110100111;
		16'b0111110011010011: color_data = 12'b001110100111;
		16'b0111110011010100: color_data = 12'b001110100111;
		16'b0111110011010101: color_data = 12'b001110100111;
		16'b0111110011010110: color_data = 12'b001110100111;
		16'b0111110011010111: color_data = 12'b001110100111;
		16'b0111110011011000: color_data = 12'b001110100111;
		16'b0111110011011001: color_data = 12'b001110100111;
		16'b0111110011011010: color_data = 12'b001110100111;
		16'b0111110011011011: color_data = 12'b001110100111;
		16'b0111110011011100: color_data = 12'b001110100111;
		16'b0111110011011101: color_data = 12'b001110100111;
		16'b0111110011011110: color_data = 12'b001110100111;
		16'b0111110011011111: color_data = 12'b001110100111;
		16'b0111110011100000: color_data = 12'b001110100111;
		16'b0111110011100001: color_data = 12'b001110100111;
		16'b0111110011100010: color_data = 12'b001110100111;
		16'b0111110011110110: color_data = 12'b001110100111;
		16'b0111110011110111: color_data = 12'b001110100111;
		16'b0111110011111000: color_data = 12'b001110100111;
		16'b0111110011111001: color_data = 12'b001110100111;
		16'b0111110011111010: color_data = 12'b001110100111;
		16'b0111110011111011: color_data = 12'b001110100111;
		16'b0111110011111100: color_data = 12'b001110100111;
		16'b0111110011111101: color_data = 12'b001110100111;
		16'b0111110011111110: color_data = 12'b001110100111;
		16'b0111110011111111: color_data = 12'b001110100111;
		16'b0111110100000000: color_data = 12'b001110100111;
		16'b0111110100000001: color_data = 12'b001110100111;
		16'b0111110100011010: color_data = 12'b001110100111;
		16'b0111110100011011: color_data = 12'b001110100111;
		16'b0111110100011100: color_data = 12'b001110100111;
		16'b0111110100011101: color_data = 12'b001110100111;
		16'b0111110100011110: color_data = 12'b001110100111;
		16'b0111110100011111: color_data = 12'b001110100111;
		16'b0111110100100000: color_data = 12'b001110100111;
		16'b0111110100100001: color_data = 12'b001110100111;
		16'b0111110100100010: color_data = 12'b001110100111;
		16'b0111110100100011: color_data = 12'b001110100111;
		16'b0111110100100100: color_data = 12'b001110100111;
		16'b0111110100100101: color_data = 12'b001110100111;
		16'b0111110100100110: color_data = 12'b001110100111;
		16'b0111110100101101: color_data = 12'b001110100111;
		16'b0111110100101110: color_data = 12'b001110100111;
		16'b0111110100101111: color_data = 12'b001110100111;
		16'b0111110100110000: color_data = 12'b001110100111;
		16'b0111110100110001: color_data = 12'b001110100111;
		16'b0111110100110010: color_data = 12'b001110100111;
		16'b0111110100110011: color_data = 12'b001110100111;
		16'b0111110100110100: color_data = 12'b001110100111;
		16'b0111110100110101: color_data = 12'b001110100111;
		16'b0111110100110110: color_data = 12'b001110100111;
		16'b0111110100110111: color_data = 12'b001110100111;
		16'b0111110100111000: color_data = 12'b001110100111;
		16'b0111110101000101: color_data = 12'b001110100111;
		16'b0111110101000110: color_data = 12'b001110100111;
		16'b0111110101000111: color_data = 12'b001110100111;
		16'b0111110101001000: color_data = 12'b001110100111;
		16'b0111110101001001: color_data = 12'b001110100111;
		16'b0111110101001010: color_data = 12'b001110100111;
		16'b0111110101001011: color_data = 12'b001110100111;
		16'b0111110101001100: color_data = 12'b001110100111;
		16'b0111110101001101: color_data = 12'b001110100111;
		16'b0111110101001110: color_data = 12'b001110100111;
		16'b0111110101001111: color_data = 12'b001110100111;
		16'b0111110101010000: color_data = 12'b001110100111;
		16'b0111110101010001: color_data = 12'b001110100111;
		16'b0111110101011000: color_data = 12'b001110100111;
		16'b0111110101011001: color_data = 12'b001110100111;
		16'b0111110101011010: color_data = 12'b001110100111;
		16'b0111110101011011: color_data = 12'b001110100111;
		16'b0111110101011100: color_data = 12'b001110100111;
		16'b0111110101011101: color_data = 12'b001110100111;
		16'b0111110101011110: color_data = 12'b001110100111;
		16'b0111110101011111: color_data = 12'b001110100111;
		16'b0111110101100000: color_data = 12'b001110100111;
		16'b0111110101100001: color_data = 12'b001110100111;
		16'b0111110101100010: color_data = 12'b001110100111;
		16'b0111110101100011: color_data = 12'b001110100111;
		16'b0111110101110000: color_data = 12'b001110100111;
		16'b0111110101110001: color_data = 12'b001110100111;
		16'b0111110101110010: color_data = 12'b001110100111;
		16'b0111110101110011: color_data = 12'b001110100111;
		16'b0111110101110100: color_data = 12'b001110100111;
		16'b0111110101110101: color_data = 12'b001110100111;
		16'b0111110101110110: color_data = 12'b001110100111;
		16'b0111110101110111: color_data = 12'b001110100111;
		16'b0111110101111000: color_data = 12'b001110100111;
		16'b0111110101111001: color_data = 12'b001110100111;
		16'b0111110101111010: color_data = 12'b001110100111;
		16'b0111110101111011: color_data = 12'b001110100111;
		16'b0111111000000000: color_data = 12'b001110100111;
		16'b0111111000000001: color_data = 12'b001110100111;
		16'b0111111000000010: color_data = 12'b001110100111;
		16'b0111111000000011: color_data = 12'b001110100111;
		16'b0111111000000100: color_data = 12'b001110100111;
		16'b0111111000000101: color_data = 12'b001110100111;
		16'b0111111000000110: color_data = 12'b001110100111;
		16'b0111111000000111: color_data = 12'b001110100111;
		16'b0111111000001000: color_data = 12'b001110100111;
		16'b0111111000001001: color_data = 12'b001110100111;
		16'b0111111000001010: color_data = 12'b001110100111;
		16'b0111111000001011: color_data = 12'b001110100111;
		16'b0111111000001100: color_data = 12'b001110100111;
		16'b0111111000101011: color_data = 12'b001110100111;
		16'b0111111000101100: color_data = 12'b001110100111;
		16'b0111111000101101: color_data = 12'b001110100111;
		16'b0111111000101110: color_data = 12'b001110100111;
		16'b0111111000101111: color_data = 12'b001110100111;
		16'b0111111000110000: color_data = 12'b001110100111;
		16'b0111111000110001: color_data = 12'b001110100111;
		16'b0111111000110010: color_data = 12'b001110100111;
		16'b0111111000110011: color_data = 12'b001110100111;
		16'b0111111000110100: color_data = 12'b001110100111;
		16'b0111111000110101: color_data = 12'b001110100111;
		16'b0111111000110110: color_data = 12'b001110100111;
		16'b0111111000110111: color_data = 12'b001110100111;
		16'b0111111000111000: color_data = 12'b001110100111;
		16'b0111111000111001: color_data = 12'b001110100111;
		16'b0111111000111010: color_data = 12'b001110100111;
		16'b0111111000111011: color_data = 12'b001110100111;
		16'b0111111000111100: color_data = 12'b001110100111;
		16'b0111111000111101: color_data = 12'b001110100111;
		16'b0111111000111110: color_data = 12'b001110100111;
		16'b0111111000111111: color_data = 12'b001110100111;
		16'b0111111001000000: color_data = 12'b001110100111;
		16'b0111111001000001: color_data = 12'b001110100111;
		16'b0111111001000010: color_data = 12'b001110100111;
		16'b0111111001000011: color_data = 12'b001110100111;
		16'b0111111001000100: color_data = 12'b001110100111;
		16'b0111111001000101: color_data = 12'b001110100111;
		16'b0111111001000110: color_data = 12'b001110100111;
		16'b0111111001000111: color_data = 12'b001110100111;
		16'b0111111001001000: color_data = 12'b001110100111;
		16'b0111111001001001: color_data = 12'b001110100111;
		16'b0111111001001010: color_data = 12'b001110100111;
		16'b0111111001001011: color_data = 12'b001110100111;
		16'b0111111001001100: color_data = 12'b001110100111;
		16'b0111111001001101: color_data = 12'b001110100111;
		16'b0111111001001110: color_data = 12'b001110100111;
		16'b0111111001001111: color_data = 12'b001110100111;
		16'b0111111001011100: color_data = 12'b001110100111;
		16'b0111111001011101: color_data = 12'b001110100111;
		16'b0111111001011110: color_data = 12'b001110100111;
		16'b0111111001011111: color_data = 12'b001110100111;
		16'b0111111001100000: color_data = 12'b001110100111;
		16'b0111111001100001: color_data = 12'b001110100111;
		16'b0111111001100010: color_data = 12'b001110100111;
		16'b0111111001100011: color_data = 12'b001110100111;
		16'b0111111001100100: color_data = 12'b001110100111;
		16'b0111111001100101: color_data = 12'b001110100111;
		16'b0111111001100110: color_data = 12'b001110100111;
		16'b0111111001100111: color_data = 12'b001110100111;
		16'b0111111001101000: color_data = 12'b001110100111;
		16'b0111111001110101: color_data = 12'b001110100111;
		16'b0111111001110110: color_data = 12'b001110100111;
		16'b0111111001110111: color_data = 12'b001110100111;
		16'b0111111001111000: color_data = 12'b001110100111;
		16'b0111111001111001: color_data = 12'b001110100111;
		16'b0111111001111010: color_data = 12'b001110100111;
		16'b0111111001111011: color_data = 12'b001110100111;
		16'b0111111001111100: color_data = 12'b001110100111;
		16'b0111111001111101: color_data = 12'b001110100111;
		16'b0111111001111110: color_data = 12'b001110100111;
		16'b0111111001111111: color_data = 12'b001110100111;
		16'b0111111010000000: color_data = 12'b001110100111;
		16'b0111111010001101: color_data = 12'b001110100111;
		16'b0111111010001110: color_data = 12'b001110100111;
		16'b0111111010001111: color_data = 12'b001110100111;
		16'b0111111010010000: color_data = 12'b001110100111;
		16'b0111111010010001: color_data = 12'b001110100111;
		16'b0111111010010010: color_data = 12'b001110100111;
		16'b0111111010010011: color_data = 12'b001110100111;
		16'b0111111010010100: color_data = 12'b001110100111;
		16'b0111111010010101: color_data = 12'b001110100111;
		16'b0111111010010110: color_data = 12'b001110100111;
		16'b0111111010010111: color_data = 12'b001110100111;
		16'b0111111010011000: color_data = 12'b001110100111;
		16'b0111111010011001: color_data = 12'b001110100111;
		16'b0111111010100000: color_data = 12'b001110100111;
		16'b0111111010100001: color_data = 12'b001110100111;
		16'b0111111010100010: color_data = 12'b001110100111;
		16'b0111111010100011: color_data = 12'b001110100111;
		16'b0111111010100100: color_data = 12'b001110100111;
		16'b0111111010100101: color_data = 12'b001110100111;
		16'b0111111010100110: color_data = 12'b001110100111;
		16'b0111111010100111: color_data = 12'b001110100111;
		16'b0111111010101000: color_data = 12'b001110100111;
		16'b0111111010101001: color_data = 12'b001110100111;
		16'b0111111010101010: color_data = 12'b001110100111;
		16'b0111111010101011: color_data = 12'b001110100111;
		16'b0111111010111000: color_data = 12'b001110100111;
		16'b0111111010111001: color_data = 12'b001110100111;
		16'b0111111010111010: color_data = 12'b001110100111;
		16'b0111111010111011: color_data = 12'b001110100111;
		16'b0111111010111100: color_data = 12'b001110100111;
		16'b0111111010111101: color_data = 12'b001110100111;
		16'b0111111010111110: color_data = 12'b001110100111;
		16'b0111111010111111: color_data = 12'b001110100111;
		16'b0111111011000000: color_data = 12'b001110100111;
		16'b0111111011000001: color_data = 12'b001110100111;
		16'b0111111011000010: color_data = 12'b001110100111;
		16'b0111111011000011: color_data = 12'b001110100111;
		16'b0111111011000100: color_data = 12'b001110100111;
		16'b0111111011001011: color_data = 12'b001110100111;
		16'b0111111011001100: color_data = 12'b001110100111;
		16'b0111111011001101: color_data = 12'b001110100111;
		16'b0111111011001110: color_data = 12'b001110100111;
		16'b0111111011001111: color_data = 12'b001110100111;
		16'b0111111011010000: color_data = 12'b001110100111;
		16'b0111111011010001: color_data = 12'b001110100111;
		16'b0111111011010010: color_data = 12'b001110100111;
		16'b0111111011010011: color_data = 12'b001110100111;
		16'b0111111011010100: color_data = 12'b001110100111;
		16'b0111111011010101: color_data = 12'b001110100111;
		16'b0111111011010110: color_data = 12'b001110100111;
		16'b0111111011010111: color_data = 12'b001110100111;
		16'b0111111011011000: color_data = 12'b001110100111;
		16'b0111111011011001: color_data = 12'b001110100111;
		16'b0111111011011010: color_data = 12'b001110100111;
		16'b0111111011011011: color_data = 12'b001110100111;
		16'b0111111011011100: color_data = 12'b001110100111;
		16'b0111111011011101: color_data = 12'b001110100111;
		16'b0111111011011110: color_data = 12'b001110100111;
		16'b0111111011011111: color_data = 12'b001110100111;
		16'b0111111011100000: color_data = 12'b001110100111;
		16'b0111111011100001: color_data = 12'b001110100111;
		16'b0111111011100010: color_data = 12'b001110100111;
		16'b0111111011110110: color_data = 12'b001110100111;
		16'b0111111011110111: color_data = 12'b001110100111;
		16'b0111111011111000: color_data = 12'b001110100111;
		16'b0111111011111001: color_data = 12'b001110100111;
		16'b0111111011111010: color_data = 12'b001110100111;
		16'b0111111011111011: color_data = 12'b001110100111;
		16'b0111111011111100: color_data = 12'b001110100111;
		16'b0111111011111101: color_data = 12'b001110100111;
		16'b0111111011111110: color_data = 12'b001110100111;
		16'b0111111011111111: color_data = 12'b001110100111;
		16'b0111111100000000: color_data = 12'b001110100111;
		16'b0111111100000001: color_data = 12'b001110100111;
		16'b0111111100011010: color_data = 12'b001110100111;
		16'b0111111100011011: color_data = 12'b001110100111;
		16'b0111111100011100: color_data = 12'b001110100111;
		16'b0111111100011101: color_data = 12'b001110100111;
		16'b0111111100011110: color_data = 12'b001110100111;
		16'b0111111100011111: color_data = 12'b001110100111;
		16'b0111111100100000: color_data = 12'b001110100111;
		16'b0111111100100001: color_data = 12'b001110100111;
		16'b0111111100100010: color_data = 12'b001110100111;
		16'b0111111100100011: color_data = 12'b001110100111;
		16'b0111111100100100: color_data = 12'b001110100111;
		16'b0111111100100101: color_data = 12'b001110100111;
		16'b0111111100100110: color_data = 12'b001110100111;
		16'b0111111100101101: color_data = 12'b001110100111;
		16'b0111111100101110: color_data = 12'b001110100111;
		16'b0111111100101111: color_data = 12'b001110100111;
		16'b0111111100110000: color_data = 12'b001110100111;
		16'b0111111100110001: color_data = 12'b001110100111;
		16'b0111111100110010: color_data = 12'b001110100111;
		16'b0111111100110011: color_data = 12'b001110100111;
		16'b0111111100110100: color_data = 12'b001110100111;
		16'b0111111100110101: color_data = 12'b001110100111;
		16'b0111111100110110: color_data = 12'b001110100111;
		16'b0111111100110111: color_data = 12'b001110100111;
		16'b0111111100111000: color_data = 12'b001110100111;
		16'b0111111101000101: color_data = 12'b001110100111;
		16'b0111111101000110: color_data = 12'b001110100111;
		16'b0111111101000111: color_data = 12'b001110100111;
		16'b0111111101001000: color_data = 12'b001110100111;
		16'b0111111101001001: color_data = 12'b001110100111;
		16'b0111111101001010: color_data = 12'b001110100111;
		16'b0111111101001011: color_data = 12'b001110100111;
		16'b0111111101001100: color_data = 12'b001110100111;
		16'b0111111101001101: color_data = 12'b001110100111;
		16'b0111111101001110: color_data = 12'b001110100111;
		16'b0111111101001111: color_data = 12'b001110100111;
		16'b0111111101010000: color_data = 12'b001110100111;
		16'b0111111101010001: color_data = 12'b001110100111;
		16'b0111111101011000: color_data = 12'b001110100111;
		16'b0111111101011001: color_data = 12'b001110100111;
		16'b0111111101011010: color_data = 12'b001110100111;
		16'b0111111101011011: color_data = 12'b001110100111;
		16'b0111111101011100: color_data = 12'b001110100111;
		16'b0111111101011101: color_data = 12'b001110100111;
		16'b0111111101011110: color_data = 12'b001110100111;
		16'b0111111101011111: color_data = 12'b001110100111;
		16'b0111111101100000: color_data = 12'b001110100111;
		16'b0111111101100001: color_data = 12'b001110100111;
		16'b0111111101100010: color_data = 12'b001110100111;
		16'b0111111101100011: color_data = 12'b001110100111;
		16'b0111111101110000: color_data = 12'b001110100111;
		16'b0111111101110001: color_data = 12'b001110100111;
		16'b0111111101110010: color_data = 12'b001110100111;
		16'b0111111101110011: color_data = 12'b001110100111;
		16'b0111111101110100: color_data = 12'b001110100111;
		16'b0111111101110101: color_data = 12'b001110100111;
		16'b0111111101110110: color_data = 12'b001110100111;
		16'b0111111101110111: color_data = 12'b001110100111;
		16'b0111111101111000: color_data = 12'b001110100111;
		16'b0111111101111001: color_data = 12'b001110100111;
		16'b0111111101111010: color_data = 12'b001110100111;
		16'b0111111101111011: color_data = 12'b001110100111;
		16'b1000000000000000: color_data = 12'b001110100111;
		16'b1000000000000001: color_data = 12'b001110100111;
		16'b1000000000000010: color_data = 12'b001110100111;
		16'b1000000000000011: color_data = 12'b001110100111;
		16'b1000000000000100: color_data = 12'b001110100111;
		16'b1000000000000101: color_data = 12'b001110100111;
		16'b1000000000000110: color_data = 12'b001110100111;
		16'b1000000000000111: color_data = 12'b001110100111;
		16'b1000000000001000: color_data = 12'b001110100111;
		16'b1000000000001001: color_data = 12'b001110100111;
		16'b1000000000001010: color_data = 12'b001110100111;
		16'b1000000000001011: color_data = 12'b001110100111;
		16'b1000000000001100: color_data = 12'b001110100111;
		16'b1000000000101011: color_data = 12'b001110100111;
		16'b1000000000101100: color_data = 12'b001110100111;
		16'b1000000000101101: color_data = 12'b001110100111;
		16'b1000000000101110: color_data = 12'b001110100111;
		16'b1000000000101111: color_data = 12'b001110100111;
		16'b1000000000110000: color_data = 12'b001110100111;
		16'b1000000000110001: color_data = 12'b001110100111;
		16'b1000000000110010: color_data = 12'b001110100111;
		16'b1000000000110011: color_data = 12'b001110100111;
		16'b1000000000110100: color_data = 12'b001110100111;
		16'b1000000000110101: color_data = 12'b001110100111;
		16'b1000000000110110: color_data = 12'b001110100111;
		16'b1000000000110111: color_data = 12'b001110100111;
		16'b1000000001000100: color_data = 12'b001110100111;
		16'b1000000001000101: color_data = 12'b001110100111;
		16'b1000000001000110: color_data = 12'b001110100111;
		16'b1000000001000111: color_data = 12'b001110100111;
		16'b1000000001001000: color_data = 12'b001110100111;
		16'b1000000001001001: color_data = 12'b001110100111;
		16'b1000000001001010: color_data = 12'b001110100111;
		16'b1000000001001011: color_data = 12'b001110100111;
		16'b1000000001001100: color_data = 12'b001110100111;
		16'b1000000001001101: color_data = 12'b001110100111;
		16'b1000000001001110: color_data = 12'b001110100111;
		16'b1000000001001111: color_data = 12'b001110100111;
		16'b1000000001011100: color_data = 12'b001110100111;
		16'b1000000001011101: color_data = 12'b001110100111;
		16'b1000000001011110: color_data = 12'b001110100111;
		16'b1000000001011111: color_data = 12'b001110100111;
		16'b1000000001100000: color_data = 12'b001110100111;
		16'b1000000001100001: color_data = 12'b001110100111;
		16'b1000000001100010: color_data = 12'b001110100111;
		16'b1000000001100011: color_data = 12'b001110100111;
		16'b1000000001100100: color_data = 12'b001110100111;
		16'b1000000001100101: color_data = 12'b001110100111;
		16'b1000000001100110: color_data = 12'b001110100111;
		16'b1000000001100111: color_data = 12'b001110100111;
		16'b1000000001101000: color_data = 12'b001110100111;
		16'b1000000001110101: color_data = 12'b001110100111;
		16'b1000000001110110: color_data = 12'b001110100111;
		16'b1000000001110111: color_data = 12'b001110100111;
		16'b1000000001111000: color_data = 12'b001110100111;
		16'b1000000001111001: color_data = 12'b001110100111;
		16'b1000000001111010: color_data = 12'b001110100111;
		16'b1000000001111011: color_data = 12'b001110100111;
		16'b1000000001111100: color_data = 12'b001110100111;
		16'b1000000001111101: color_data = 12'b001110100111;
		16'b1000000001111110: color_data = 12'b001110100111;
		16'b1000000001111111: color_data = 12'b001110100111;
		16'b1000000010000000: color_data = 12'b001110100111;
		16'b1000000010001101: color_data = 12'b001110100111;
		16'b1000000010001110: color_data = 12'b001110100111;
		16'b1000000010001111: color_data = 12'b001110100111;
		16'b1000000010010000: color_data = 12'b001110100111;
		16'b1000000010010001: color_data = 12'b001110100111;
		16'b1000000010010010: color_data = 12'b001110100111;
		16'b1000000010010011: color_data = 12'b001110100111;
		16'b1000000010010100: color_data = 12'b001110100111;
		16'b1000000010010101: color_data = 12'b001110100111;
		16'b1000000010010110: color_data = 12'b001110100111;
		16'b1000000010010111: color_data = 12'b001110100111;
		16'b1000000010011000: color_data = 12'b001110100111;
		16'b1000000010011001: color_data = 12'b001110100111;
		16'b1000000010100000: color_data = 12'b001110100111;
		16'b1000000010100001: color_data = 12'b001110100111;
		16'b1000000010100010: color_data = 12'b001110100111;
		16'b1000000010100011: color_data = 12'b001110100111;
		16'b1000000010100100: color_data = 12'b001110100111;
		16'b1000000010100101: color_data = 12'b001110100111;
		16'b1000000010100110: color_data = 12'b001110100111;
		16'b1000000010100111: color_data = 12'b001110100111;
		16'b1000000010101000: color_data = 12'b001110100111;
		16'b1000000010101001: color_data = 12'b001110100111;
		16'b1000000010101010: color_data = 12'b001110100111;
		16'b1000000010101011: color_data = 12'b001110100111;
		16'b1000000010111000: color_data = 12'b001110100111;
		16'b1000000010111001: color_data = 12'b001110100111;
		16'b1000000010111010: color_data = 12'b001110100111;
		16'b1000000010111011: color_data = 12'b001110100111;
		16'b1000000010111100: color_data = 12'b001110100111;
		16'b1000000010111101: color_data = 12'b001110100111;
		16'b1000000010111110: color_data = 12'b001110100111;
		16'b1000000010111111: color_data = 12'b001110100111;
		16'b1000000011000000: color_data = 12'b001110100111;
		16'b1000000011000001: color_data = 12'b001110100111;
		16'b1000000011000010: color_data = 12'b001110100111;
		16'b1000000011000011: color_data = 12'b001110100111;
		16'b1000000011000100: color_data = 12'b001110100111;
		16'b1000000011001011: color_data = 12'b001110100111;
		16'b1000000011001100: color_data = 12'b001110100111;
		16'b1000000011001101: color_data = 12'b001110100111;
		16'b1000000011001110: color_data = 12'b001110100111;
		16'b1000000011001111: color_data = 12'b001110100111;
		16'b1000000011010000: color_data = 12'b001110100111;
		16'b1000000011010001: color_data = 12'b001110100111;
		16'b1000000011010010: color_data = 12'b001110100111;
		16'b1000000011010011: color_data = 12'b001110100111;
		16'b1000000011010100: color_data = 12'b001110100111;
		16'b1000000011010101: color_data = 12'b001110100111;
		16'b1000000011010110: color_data = 12'b001110100111;
		16'b1000000011110110: color_data = 12'b001110100111;
		16'b1000000011110111: color_data = 12'b001110100111;
		16'b1000000011111000: color_data = 12'b001110100111;
		16'b1000000011111001: color_data = 12'b001110100111;
		16'b1000000011111010: color_data = 12'b001110100111;
		16'b1000000011111011: color_data = 12'b001110100111;
		16'b1000000011111100: color_data = 12'b001110100111;
		16'b1000000011111101: color_data = 12'b001110100111;
		16'b1000000011111110: color_data = 12'b001110100111;
		16'b1000000011111111: color_data = 12'b001110100111;
		16'b1000000100000000: color_data = 12'b001110100111;
		16'b1000000100000001: color_data = 12'b001110100111;
		16'b1000000100011010: color_data = 12'b001110100111;
		16'b1000000100011011: color_data = 12'b001110100111;
		16'b1000000100011100: color_data = 12'b001110100111;
		16'b1000000100011101: color_data = 12'b001110100111;
		16'b1000000100011110: color_data = 12'b001110100111;
		16'b1000000100011111: color_data = 12'b001110100111;
		16'b1000000100100000: color_data = 12'b001110100111;
		16'b1000000100100001: color_data = 12'b001110100111;
		16'b1000000100100010: color_data = 12'b001110100111;
		16'b1000000100100011: color_data = 12'b001110100111;
		16'b1000000100100100: color_data = 12'b001110100111;
		16'b1000000100100101: color_data = 12'b001110100111;
		16'b1000000100100110: color_data = 12'b001110100111;
		16'b1000000100101101: color_data = 12'b001110100111;
		16'b1000000100101110: color_data = 12'b001110100111;
		16'b1000000100101111: color_data = 12'b001110100111;
		16'b1000000100110000: color_data = 12'b001110100111;
		16'b1000000100110001: color_data = 12'b001110100111;
		16'b1000000100110010: color_data = 12'b001110100111;
		16'b1000000100110011: color_data = 12'b001110100111;
		16'b1000000100110100: color_data = 12'b001110100111;
		16'b1000000100110101: color_data = 12'b001110100111;
		16'b1000000100110110: color_data = 12'b001110100111;
		16'b1000000100110111: color_data = 12'b001110100111;
		16'b1000000100111000: color_data = 12'b001110100111;
		16'b1000000101000101: color_data = 12'b001110100111;
		16'b1000000101000110: color_data = 12'b001110100111;
		16'b1000000101000111: color_data = 12'b001110100111;
		16'b1000000101001000: color_data = 12'b001110100111;
		16'b1000000101001001: color_data = 12'b001110100111;
		16'b1000000101001010: color_data = 12'b001110100111;
		16'b1000000101001011: color_data = 12'b001110100111;
		16'b1000000101001100: color_data = 12'b001110100111;
		16'b1000000101001101: color_data = 12'b001110100111;
		16'b1000000101001110: color_data = 12'b001110100111;
		16'b1000000101001111: color_data = 12'b001110100111;
		16'b1000000101010000: color_data = 12'b001110100111;
		16'b1000000101010001: color_data = 12'b001110100111;
		16'b1000000101011000: color_data = 12'b001110100111;
		16'b1000000101011001: color_data = 12'b001110100111;
		16'b1000000101011010: color_data = 12'b001110100111;
		16'b1000000101011011: color_data = 12'b001110100111;
		16'b1000000101011100: color_data = 12'b001110100111;
		16'b1000000101011101: color_data = 12'b001110100111;
		16'b1000000101011110: color_data = 12'b001110100111;
		16'b1000000101011111: color_data = 12'b001110100111;
		16'b1000000101100000: color_data = 12'b001110100111;
		16'b1000000101100001: color_data = 12'b001110100111;
		16'b1000000101100010: color_data = 12'b001110100111;
		16'b1000000101100011: color_data = 12'b001110100111;
		16'b1000000101110000: color_data = 12'b001110100111;
		16'b1000000101110001: color_data = 12'b001110100111;
		16'b1000000101110010: color_data = 12'b001110100111;
		16'b1000000101110011: color_data = 12'b001110100111;
		16'b1000000101110100: color_data = 12'b001110100111;
		16'b1000000101110101: color_data = 12'b001110100111;
		16'b1000000101110110: color_data = 12'b001110100111;
		16'b1000000101110111: color_data = 12'b001110100111;
		16'b1000000101111000: color_data = 12'b001110100111;
		16'b1000000101111001: color_data = 12'b001110100111;
		16'b1000000101111010: color_data = 12'b001110100111;
		16'b1000000101111011: color_data = 12'b001110100111;
		16'b1000001000000000: color_data = 12'b001110100111;
		16'b1000001000000001: color_data = 12'b001110100111;
		16'b1000001000000010: color_data = 12'b001110100111;
		16'b1000001000000011: color_data = 12'b001110100111;
		16'b1000001000000100: color_data = 12'b001110100111;
		16'b1000001000000101: color_data = 12'b001110100111;
		16'b1000001000000110: color_data = 12'b001110100111;
		16'b1000001000000111: color_data = 12'b001110100111;
		16'b1000001000001000: color_data = 12'b001110100111;
		16'b1000001000001001: color_data = 12'b001110100111;
		16'b1000001000001010: color_data = 12'b001110100111;
		16'b1000001000001011: color_data = 12'b001110100111;
		16'b1000001000001100: color_data = 12'b001110100111;
		16'b1000001000101011: color_data = 12'b001110100111;
		16'b1000001000101100: color_data = 12'b001110100111;
		16'b1000001000101101: color_data = 12'b001110100111;
		16'b1000001000101110: color_data = 12'b001110100111;
		16'b1000001000101111: color_data = 12'b001110100111;
		16'b1000001000110000: color_data = 12'b001110100111;
		16'b1000001000110001: color_data = 12'b001110100111;
		16'b1000001000110010: color_data = 12'b001110100111;
		16'b1000001000110011: color_data = 12'b001110100111;
		16'b1000001000110100: color_data = 12'b001110100111;
		16'b1000001000110101: color_data = 12'b001110100111;
		16'b1000001000110110: color_data = 12'b001110100111;
		16'b1000001000110111: color_data = 12'b001110100111;
		16'b1000001001000100: color_data = 12'b001110100111;
		16'b1000001001000101: color_data = 12'b001110100111;
		16'b1000001001000110: color_data = 12'b001110100111;
		16'b1000001001000111: color_data = 12'b001110100111;
		16'b1000001001001000: color_data = 12'b001110100111;
		16'b1000001001001001: color_data = 12'b001110100111;
		16'b1000001001001010: color_data = 12'b001110100111;
		16'b1000001001001011: color_data = 12'b001110100111;
		16'b1000001001001100: color_data = 12'b001110100111;
		16'b1000001001001101: color_data = 12'b001110100111;
		16'b1000001001001110: color_data = 12'b001110100111;
		16'b1000001001001111: color_data = 12'b001110100111;
		16'b1000001001011100: color_data = 12'b001110100111;
		16'b1000001001011101: color_data = 12'b001110100111;
		16'b1000001001011110: color_data = 12'b001110100111;
		16'b1000001001011111: color_data = 12'b001110100111;
		16'b1000001001100000: color_data = 12'b001110100111;
		16'b1000001001100001: color_data = 12'b001110100111;
		16'b1000001001100010: color_data = 12'b001110100111;
		16'b1000001001100011: color_data = 12'b001110100111;
		16'b1000001001100100: color_data = 12'b001110100111;
		16'b1000001001100101: color_data = 12'b001110100111;
		16'b1000001001100110: color_data = 12'b001110100111;
		16'b1000001001100111: color_data = 12'b001110100111;
		16'b1000001001101000: color_data = 12'b001110100111;
		16'b1000001001110101: color_data = 12'b001110100111;
		16'b1000001001110110: color_data = 12'b001110100111;
		16'b1000001001110111: color_data = 12'b001110100111;
		16'b1000001001111000: color_data = 12'b001110100111;
		16'b1000001001111001: color_data = 12'b001110100111;
		16'b1000001001111010: color_data = 12'b001110100111;
		16'b1000001001111011: color_data = 12'b001110100111;
		16'b1000001001111100: color_data = 12'b001110100111;
		16'b1000001001111101: color_data = 12'b001110100111;
		16'b1000001001111110: color_data = 12'b001110100111;
		16'b1000001001111111: color_data = 12'b001110100111;
		16'b1000001010000000: color_data = 12'b001110100111;
		16'b1000001010001101: color_data = 12'b001110100111;
		16'b1000001010001110: color_data = 12'b001110100111;
		16'b1000001010001111: color_data = 12'b001110100111;
		16'b1000001010010000: color_data = 12'b001110100111;
		16'b1000001010010001: color_data = 12'b001110100111;
		16'b1000001010010010: color_data = 12'b001110100111;
		16'b1000001010010011: color_data = 12'b001110100111;
		16'b1000001010010100: color_data = 12'b001110100111;
		16'b1000001010010101: color_data = 12'b001110100111;
		16'b1000001010010110: color_data = 12'b001110100111;
		16'b1000001010010111: color_data = 12'b001110100111;
		16'b1000001010011000: color_data = 12'b001110100111;
		16'b1000001010011001: color_data = 12'b001110100111;
		16'b1000001010100000: color_data = 12'b001110100111;
		16'b1000001010100001: color_data = 12'b001110100111;
		16'b1000001010100010: color_data = 12'b001110100111;
		16'b1000001010100011: color_data = 12'b001110100111;
		16'b1000001010100100: color_data = 12'b001110100111;
		16'b1000001010100101: color_data = 12'b001110100111;
		16'b1000001010100110: color_data = 12'b001110100111;
		16'b1000001010100111: color_data = 12'b001110100111;
		16'b1000001010101000: color_data = 12'b001110100111;
		16'b1000001010101001: color_data = 12'b001110100111;
		16'b1000001010101010: color_data = 12'b001110100111;
		16'b1000001010101011: color_data = 12'b001110100111;
		16'b1000001010111000: color_data = 12'b001110100111;
		16'b1000001010111001: color_data = 12'b001110100111;
		16'b1000001010111010: color_data = 12'b001110100111;
		16'b1000001010111011: color_data = 12'b001110100111;
		16'b1000001010111100: color_data = 12'b001110100111;
		16'b1000001010111101: color_data = 12'b001110100111;
		16'b1000001010111110: color_data = 12'b001110100111;
		16'b1000001010111111: color_data = 12'b001110100111;
		16'b1000001011000000: color_data = 12'b001110100111;
		16'b1000001011000001: color_data = 12'b001110100111;
		16'b1000001011000010: color_data = 12'b001110100111;
		16'b1000001011000011: color_data = 12'b001110100111;
		16'b1000001011000100: color_data = 12'b001110100111;
		16'b1000001011001011: color_data = 12'b001110100111;
		16'b1000001011001100: color_data = 12'b001110100111;
		16'b1000001011001101: color_data = 12'b001110100111;
		16'b1000001011001110: color_data = 12'b001110100111;
		16'b1000001011001111: color_data = 12'b001110100111;
		16'b1000001011010000: color_data = 12'b001110100111;
		16'b1000001011010001: color_data = 12'b001110100111;
		16'b1000001011010010: color_data = 12'b001110100111;
		16'b1000001011010011: color_data = 12'b001110100111;
		16'b1000001011010100: color_data = 12'b001110100111;
		16'b1000001011010101: color_data = 12'b001110100111;
		16'b1000001011010110: color_data = 12'b001110100111;
		16'b1000001011110110: color_data = 12'b001110100111;
		16'b1000001011110111: color_data = 12'b001110100111;
		16'b1000001011111000: color_data = 12'b001110100111;
		16'b1000001011111001: color_data = 12'b001110100111;
		16'b1000001011111010: color_data = 12'b001110100111;
		16'b1000001011111011: color_data = 12'b001110100111;
		16'b1000001011111100: color_data = 12'b001110100111;
		16'b1000001011111101: color_data = 12'b001110100111;
		16'b1000001011111110: color_data = 12'b001110100111;
		16'b1000001011111111: color_data = 12'b001110100111;
		16'b1000001100000000: color_data = 12'b001110100111;
		16'b1000001100000001: color_data = 12'b001110100111;
		16'b1000001100011010: color_data = 12'b001110100111;
		16'b1000001100011011: color_data = 12'b001110100111;
		16'b1000001100011100: color_data = 12'b001110100111;
		16'b1000001100011101: color_data = 12'b001110100111;
		16'b1000001100011110: color_data = 12'b001110100111;
		16'b1000001100011111: color_data = 12'b001110100111;
		16'b1000001100100000: color_data = 12'b001110100111;
		16'b1000001100100001: color_data = 12'b001110100111;
		16'b1000001100100010: color_data = 12'b001110100111;
		16'b1000001100100011: color_data = 12'b001110100111;
		16'b1000001100100100: color_data = 12'b001110100111;
		16'b1000001100100101: color_data = 12'b001110100111;
		16'b1000001100100110: color_data = 12'b001110100111;
		16'b1000001100101101: color_data = 12'b001110100111;
		16'b1000001100101110: color_data = 12'b001110100111;
		16'b1000001100101111: color_data = 12'b001110100111;
		16'b1000001100110000: color_data = 12'b001110100111;
		16'b1000001100110001: color_data = 12'b001110100111;
		16'b1000001100110010: color_data = 12'b001110100111;
		16'b1000001100110011: color_data = 12'b001110100111;
		16'b1000001100110100: color_data = 12'b001110100111;
		16'b1000001100110101: color_data = 12'b001110100111;
		16'b1000001100110110: color_data = 12'b001110100111;
		16'b1000001100110111: color_data = 12'b001110100111;
		16'b1000001100111000: color_data = 12'b001110100111;
		16'b1000001101000101: color_data = 12'b001110100111;
		16'b1000001101000110: color_data = 12'b001110100111;
		16'b1000001101000111: color_data = 12'b001110100111;
		16'b1000001101001000: color_data = 12'b001110100111;
		16'b1000001101001001: color_data = 12'b001110100111;
		16'b1000001101001010: color_data = 12'b001110100111;
		16'b1000001101001011: color_data = 12'b001110100111;
		16'b1000001101001100: color_data = 12'b001110100111;
		16'b1000001101001101: color_data = 12'b001110100111;
		16'b1000001101001110: color_data = 12'b001110100111;
		16'b1000001101001111: color_data = 12'b001110100111;
		16'b1000001101010000: color_data = 12'b001110100111;
		16'b1000001101010001: color_data = 12'b001110100111;
		16'b1000001101011000: color_data = 12'b001110100111;
		16'b1000001101011001: color_data = 12'b001110100111;
		16'b1000001101011010: color_data = 12'b001110100111;
		16'b1000001101011011: color_data = 12'b001110100111;
		16'b1000001101011100: color_data = 12'b001110100111;
		16'b1000001101011101: color_data = 12'b001110100111;
		16'b1000001101011110: color_data = 12'b001110100111;
		16'b1000001101011111: color_data = 12'b001110100111;
		16'b1000001101100000: color_data = 12'b001110100111;
		16'b1000001101100001: color_data = 12'b001110100111;
		16'b1000001101100010: color_data = 12'b001110100111;
		16'b1000001101100011: color_data = 12'b001110100111;
		16'b1000001101110000: color_data = 12'b001110100111;
		16'b1000001101110001: color_data = 12'b001110100111;
		16'b1000001101110010: color_data = 12'b001110100111;
		16'b1000001101110011: color_data = 12'b001110100111;
		16'b1000001101110100: color_data = 12'b001110100111;
		16'b1000001101110101: color_data = 12'b001110100111;
		16'b1000001101110110: color_data = 12'b001110100111;
		16'b1000001101110111: color_data = 12'b001110100111;
		16'b1000001101111000: color_data = 12'b001110100111;
		16'b1000001101111001: color_data = 12'b001110100111;
		16'b1000001101111010: color_data = 12'b001110100111;
		16'b1000001101111011: color_data = 12'b001110100111;
		16'b1000010000000000: color_data = 12'b001110100111;
		16'b1000010000000001: color_data = 12'b001110100111;
		16'b1000010000000010: color_data = 12'b001110100111;
		16'b1000010000000011: color_data = 12'b001110100111;
		16'b1000010000000100: color_data = 12'b001110100111;
		16'b1000010000000101: color_data = 12'b001110100111;
		16'b1000010000000110: color_data = 12'b001110100111;
		16'b1000010000000111: color_data = 12'b001110100111;
		16'b1000010000001000: color_data = 12'b001110100111;
		16'b1000010000001001: color_data = 12'b001110100111;
		16'b1000010000001010: color_data = 12'b001110100111;
		16'b1000010000001011: color_data = 12'b001110100111;
		16'b1000010000001100: color_data = 12'b001110100111;
		16'b1000010000101011: color_data = 12'b001110100111;
		16'b1000010000101100: color_data = 12'b001110100111;
		16'b1000010000101101: color_data = 12'b001110100111;
		16'b1000010000101110: color_data = 12'b001110100111;
		16'b1000010000101111: color_data = 12'b001110100111;
		16'b1000010000110000: color_data = 12'b001110100111;
		16'b1000010000110001: color_data = 12'b001110100111;
		16'b1000010000110010: color_data = 12'b001110100111;
		16'b1000010000110011: color_data = 12'b001110100111;
		16'b1000010000110100: color_data = 12'b001110100111;
		16'b1000010000110101: color_data = 12'b001110100111;
		16'b1000010000110110: color_data = 12'b001110100111;
		16'b1000010000110111: color_data = 12'b001110100111;
		16'b1000010001000100: color_data = 12'b001110100111;
		16'b1000010001000101: color_data = 12'b001110100111;
		16'b1000010001000110: color_data = 12'b001110100111;
		16'b1000010001000111: color_data = 12'b001110100111;
		16'b1000010001001000: color_data = 12'b001110100111;
		16'b1000010001001001: color_data = 12'b001110100111;
		16'b1000010001001010: color_data = 12'b001110100111;
		16'b1000010001001011: color_data = 12'b001110100111;
		16'b1000010001001100: color_data = 12'b001110100111;
		16'b1000010001001101: color_data = 12'b001110100111;
		16'b1000010001001110: color_data = 12'b001110100111;
		16'b1000010001001111: color_data = 12'b001110100111;
		16'b1000010001011100: color_data = 12'b001110100111;
		16'b1000010001011101: color_data = 12'b001110100111;
		16'b1000010001011110: color_data = 12'b001110100111;
		16'b1000010001011111: color_data = 12'b001110100111;
		16'b1000010001100000: color_data = 12'b001110100111;
		16'b1000010001100001: color_data = 12'b001110100111;
		16'b1000010001100010: color_data = 12'b001110100111;
		16'b1000010001100011: color_data = 12'b001110100111;
		16'b1000010001100100: color_data = 12'b001110100111;
		16'b1000010001100101: color_data = 12'b001110100111;
		16'b1000010001100110: color_data = 12'b001110100111;
		16'b1000010001100111: color_data = 12'b001110100111;
		16'b1000010001101000: color_data = 12'b001110100111;
		16'b1000010001110101: color_data = 12'b001110100111;
		16'b1000010001110110: color_data = 12'b001110100111;
		16'b1000010001110111: color_data = 12'b001110100111;
		16'b1000010001111000: color_data = 12'b001110100111;
		16'b1000010001111001: color_data = 12'b001110100111;
		16'b1000010001111010: color_data = 12'b001110100111;
		16'b1000010001111011: color_data = 12'b001110100111;
		16'b1000010001111100: color_data = 12'b001110100111;
		16'b1000010001111101: color_data = 12'b001110100111;
		16'b1000010001111110: color_data = 12'b001110100111;
		16'b1000010001111111: color_data = 12'b001110100111;
		16'b1000010010000000: color_data = 12'b001110100111;
		16'b1000010010001101: color_data = 12'b001110100111;
		16'b1000010010001110: color_data = 12'b001110100111;
		16'b1000010010001111: color_data = 12'b001110100111;
		16'b1000010010010000: color_data = 12'b001110100111;
		16'b1000010010010001: color_data = 12'b001110100111;
		16'b1000010010010010: color_data = 12'b001110100111;
		16'b1000010010010011: color_data = 12'b001110100111;
		16'b1000010010010100: color_data = 12'b001110100111;
		16'b1000010010010101: color_data = 12'b001110100111;
		16'b1000010010010110: color_data = 12'b001110100111;
		16'b1000010010010111: color_data = 12'b001110100111;
		16'b1000010010011000: color_data = 12'b001110100111;
		16'b1000010010011001: color_data = 12'b001110100111;
		16'b1000010010100000: color_data = 12'b001110100111;
		16'b1000010010100001: color_data = 12'b001110100111;
		16'b1000010010100010: color_data = 12'b001110100111;
		16'b1000010010100011: color_data = 12'b001110100111;
		16'b1000010010100100: color_data = 12'b001110100111;
		16'b1000010010100101: color_data = 12'b001110100111;
		16'b1000010010100110: color_data = 12'b001110100111;
		16'b1000010010100111: color_data = 12'b001110100111;
		16'b1000010010101000: color_data = 12'b001110100111;
		16'b1000010010101001: color_data = 12'b001110100111;
		16'b1000010010101010: color_data = 12'b001110100111;
		16'b1000010010101011: color_data = 12'b001110100111;
		16'b1000010010111000: color_data = 12'b001110100111;
		16'b1000010010111001: color_data = 12'b001110100111;
		16'b1000010010111010: color_data = 12'b001110100111;
		16'b1000010010111011: color_data = 12'b001110100111;
		16'b1000010010111100: color_data = 12'b001110100111;
		16'b1000010010111101: color_data = 12'b001110100111;
		16'b1000010010111110: color_data = 12'b001110100111;
		16'b1000010010111111: color_data = 12'b001110100111;
		16'b1000010011000000: color_data = 12'b001110100111;
		16'b1000010011000001: color_data = 12'b001110100111;
		16'b1000010011000010: color_data = 12'b001110100111;
		16'b1000010011000011: color_data = 12'b001110100111;
		16'b1000010011000100: color_data = 12'b001110100111;
		16'b1000010011001011: color_data = 12'b001110100111;
		16'b1000010011001100: color_data = 12'b001110100111;
		16'b1000010011001101: color_data = 12'b001110100111;
		16'b1000010011001110: color_data = 12'b001110100111;
		16'b1000010011001111: color_data = 12'b001110100111;
		16'b1000010011010000: color_data = 12'b001110100111;
		16'b1000010011010001: color_data = 12'b001110100111;
		16'b1000010011010010: color_data = 12'b001110100111;
		16'b1000010011010011: color_data = 12'b001110100111;
		16'b1000010011010100: color_data = 12'b001110100111;
		16'b1000010011010101: color_data = 12'b001110100111;
		16'b1000010011010110: color_data = 12'b001110100111;
		16'b1000010011110110: color_data = 12'b001110100111;
		16'b1000010011110111: color_data = 12'b001110100111;
		16'b1000010011111000: color_data = 12'b001110100111;
		16'b1000010011111001: color_data = 12'b001110100111;
		16'b1000010011111010: color_data = 12'b001110100111;
		16'b1000010011111011: color_data = 12'b001110100111;
		16'b1000010011111100: color_data = 12'b001110100111;
		16'b1000010011111101: color_data = 12'b001110100111;
		16'b1000010011111110: color_data = 12'b001110100111;
		16'b1000010011111111: color_data = 12'b001110100111;
		16'b1000010100000000: color_data = 12'b001110100111;
		16'b1000010100000001: color_data = 12'b001110100111;
		16'b1000010100011010: color_data = 12'b001110100111;
		16'b1000010100011011: color_data = 12'b001110100111;
		16'b1000010100011100: color_data = 12'b001110100111;
		16'b1000010100011101: color_data = 12'b001110100111;
		16'b1000010100011110: color_data = 12'b001110100111;
		16'b1000010100011111: color_data = 12'b001110100111;
		16'b1000010100100000: color_data = 12'b001110100111;
		16'b1000010100100001: color_data = 12'b001110100111;
		16'b1000010100100010: color_data = 12'b001110100111;
		16'b1000010100100011: color_data = 12'b001110100111;
		16'b1000010100100100: color_data = 12'b001110100111;
		16'b1000010100100101: color_data = 12'b001110100111;
		16'b1000010100100110: color_data = 12'b001110100111;
		16'b1000010100101101: color_data = 12'b001110100111;
		16'b1000010100101110: color_data = 12'b001110100111;
		16'b1000010100101111: color_data = 12'b001110100111;
		16'b1000010100110000: color_data = 12'b001110100111;
		16'b1000010100110001: color_data = 12'b001110100111;
		16'b1000010100110010: color_data = 12'b001110100111;
		16'b1000010100110011: color_data = 12'b001110100111;
		16'b1000010100110100: color_data = 12'b001110100111;
		16'b1000010100110101: color_data = 12'b001110100111;
		16'b1000010100110110: color_data = 12'b001110100111;
		16'b1000010100110111: color_data = 12'b001110100111;
		16'b1000010100111000: color_data = 12'b001110100111;
		16'b1000010101000101: color_data = 12'b001110100111;
		16'b1000010101000110: color_data = 12'b001110100111;
		16'b1000010101000111: color_data = 12'b001110100111;
		16'b1000010101001000: color_data = 12'b001110100111;
		16'b1000010101001001: color_data = 12'b001110100111;
		16'b1000010101001010: color_data = 12'b001110100111;
		16'b1000010101001011: color_data = 12'b001110100111;
		16'b1000010101001100: color_data = 12'b001110100111;
		16'b1000010101001101: color_data = 12'b001110100111;
		16'b1000010101001110: color_data = 12'b001110100111;
		16'b1000010101001111: color_data = 12'b001110100111;
		16'b1000010101010000: color_data = 12'b001110100111;
		16'b1000010101010001: color_data = 12'b001110100111;
		16'b1000010101011000: color_data = 12'b001110100111;
		16'b1000010101011001: color_data = 12'b001110100111;
		16'b1000010101011010: color_data = 12'b001110100111;
		16'b1000010101011011: color_data = 12'b001110100111;
		16'b1000010101011100: color_data = 12'b001110100111;
		16'b1000010101011101: color_data = 12'b001110100111;
		16'b1000010101011110: color_data = 12'b001110100111;
		16'b1000010101011111: color_data = 12'b001110100111;
		16'b1000010101100000: color_data = 12'b001110100111;
		16'b1000010101100001: color_data = 12'b001110100111;
		16'b1000010101100010: color_data = 12'b001110100111;
		16'b1000010101100011: color_data = 12'b001110100111;
		16'b1000010101110000: color_data = 12'b001110100111;
		16'b1000010101110001: color_data = 12'b001110100111;
		16'b1000010101110010: color_data = 12'b001110100111;
		16'b1000010101110011: color_data = 12'b001110100111;
		16'b1000010101110100: color_data = 12'b001110100111;
		16'b1000010101110101: color_data = 12'b001110100111;
		16'b1000010101110110: color_data = 12'b001110100111;
		16'b1000010101110111: color_data = 12'b001110100111;
		16'b1000010101111000: color_data = 12'b001110100111;
		16'b1000010101111001: color_data = 12'b001110100111;
		16'b1000010101111010: color_data = 12'b001110100111;
		16'b1000010101111011: color_data = 12'b001110100111;
		16'b1000011000000000: color_data = 12'b001110100111;
		16'b1000011000000001: color_data = 12'b001110100111;
		16'b1000011000000010: color_data = 12'b001110100111;
		16'b1000011000000011: color_data = 12'b001110100111;
		16'b1000011000000100: color_data = 12'b001110100111;
		16'b1000011000000101: color_data = 12'b001110100111;
		16'b1000011000000110: color_data = 12'b001110100111;
		16'b1000011000000111: color_data = 12'b001110100111;
		16'b1000011000001000: color_data = 12'b001110100111;
		16'b1000011000001001: color_data = 12'b001110100111;
		16'b1000011000001010: color_data = 12'b001110100111;
		16'b1000011000001011: color_data = 12'b001110100111;
		16'b1000011000001100: color_data = 12'b001110100111;
		16'b1000011000101011: color_data = 12'b001110100111;
		16'b1000011000101100: color_data = 12'b001110100111;
		16'b1000011000101101: color_data = 12'b001110100111;
		16'b1000011000101110: color_data = 12'b001110100111;
		16'b1000011000101111: color_data = 12'b001110100111;
		16'b1000011000110000: color_data = 12'b001110100111;
		16'b1000011000110001: color_data = 12'b001110100111;
		16'b1000011000110010: color_data = 12'b001110100111;
		16'b1000011000110011: color_data = 12'b001110100111;
		16'b1000011000110100: color_data = 12'b001110100111;
		16'b1000011000110101: color_data = 12'b001110100111;
		16'b1000011000110110: color_data = 12'b001110100111;
		16'b1000011000110111: color_data = 12'b001110100111;
		16'b1000011001000100: color_data = 12'b001110100111;
		16'b1000011001000101: color_data = 12'b001110100111;
		16'b1000011001000110: color_data = 12'b001110100111;
		16'b1000011001000111: color_data = 12'b001110100111;
		16'b1000011001001000: color_data = 12'b001110100111;
		16'b1000011001001001: color_data = 12'b001110100111;
		16'b1000011001001010: color_data = 12'b001110100111;
		16'b1000011001001011: color_data = 12'b001110100111;
		16'b1000011001001100: color_data = 12'b001110100111;
		16'b1000011001001101: color_data = 12'b001110100111;
		16'b1000011001001110: color_data = 12'b001110100111;
		16'b1000011001001111: color_data = 12'b001110100111;
		16'b1000011001011100: color_data = 12'b001110100111;
		16'b1000011001011101: color_data = 12'b001110100111;
		16'b1000011001011110: color_data = 12'b001110100111;
		16'b1000011001011111: color_data = 12'b001110100111;
		16'b1000011001100000: color_data = 12'b001110100111;
		16'b1000011001100001: color_data = 12'b001110100111;
		16'b1000011001100010: color_data = 12'b001110100111;
		16'b1000011001100011: color_data = 12'b001110100111;
		16'b1000011001100100: color_data = 12'b001110100111;
		16'b1000011001100101: color_data = 12'b001110100111;
		16'b1000011001100110: color_data = 12'b001110100111;
		16'b1000011001100111: color_data = 12'b001110100111;
		16'b1000011001101000: color_data = 12'b001110100111;
		16'b1000011001110101: color_data = 12'b001110100111;
		16'b1000011001110110: color_data = 12'b001110100111;
		16'b1000011001110111: color_data = 12'b001110100111;
		16'b1000011001111000: color_data = 12'b001110100111;
		16'b1000011001111001: color_data = 12'b001110100111;
		16'b1000011001111010: color_data = 12'b001110100111;
		16'b1000011001111011: color_data = 12'b001110100111;
		16'b1000011001111100: color_data = 12'b001110100111;
		16'b1000011001111101: color_data = 12'b001110100111;
		16'b1000011001111110: color_data = 12'b001110100111;
		16'b1000011001111111: color_data = 12'b001110100111;
		16'b1000011010000000: color_data = 12'b001110100111;
		16'b1000011010001101: color_data = 12'b001110100111;
		16'b1000011010001110: color_data = 12'b001110100111;
		16'b1000011010001111: color_data = 12'b001110100111;
		16'b1000011010010000: color_data = 12'b001110100111;
		16'b1000011010010001: color_data = 12'b001110100111;
		16'b1000011010010010: color_data = 12'b001110100111;
		16'b1000011010010011: color_data = 12'b001110100111;
		16'b1000011010010100: color_data = 12'b001110100111;
		16'b1000011010010101: color_data = 12'b001110100111;
		16'b1000011010010110: color_data = 12'b001110100111;
		16'b1000011010010111: color_data = 12'b001110100111;
		16'b1000011010011000: color_data = 12'b001110100111;
		16'b1000011010011001: color_data = 12'b001110100111;
		16'b1000011010100000: color_data = 12'b001110100111;
		16'b1000011010100001: color_data = 12'b001110100111;
		16'b1000011010100010: color_data = 12'b001110100111;
		16'b1000011010100011: color_data = 12'b001110100111;
		16'b1000011010100100: color_data = 12'b001110100111;
		16'b1000011010100101: color_data = 12'b001110100111;
		16'b1000011010100110: color_data = 12'b001110100111;
		16'b1000011010100111: color_data = 12'b001110100111;
		16'b1000011010101000: color_data = 12'b001110100111;
		16'b1000011010101001: color_data = 12'b001110100111;
		16'b1000011010101010: color_data = 12'b001110100111;
		16'b1000011010101011: color_data = 12'b001110100111;
		16'b1000011010111000: color_data = 12'b001110100111;
		16'b1000011010111001: color_data = 12'b001110100111;
		16'b1000011010111010: color_data = 12'b001110100111;
		16'b1000011010111011: color_data = 12'b001110100111;
		16'b1000011010111100: color_data = 12'b001110100111;
		16'b1000011010111101: color_data = 12'b001110100111;
		16'b1000011010111110: color_data = 12'b001110100111;
		16'b1000011010111111: color_data = 12'b001110100111;
		16'b1000011011000000: color_data = 12'b001110100111;
		16'b1000011011000001: color_data = 12'b001110100111;
		16'b1000011011000010: color_data = 12'b001110100111;
		16'b1000011011000011: color_data = 12'b001110100111;
		16'b1000011011000100: color_data = 12'b001110100111;
		16'b1000011011001011: color_data = 12'b001110100111;
		16'b1000011011001100: color_data = 12'b001110100111;
		16'b1000011011001101: color_data = 12'b001110100111;
		16'b1000011011001110: color_data = 12'b001110100111;
		16'b1000011011001111: color_data = 12'b001110100111;
		16'b1000011011010000: color_data = 12'b001110100111;
		16'b1000011011010001: color_data = 12'b001110100111;
		16'b1000011011010010: color_data = 12'b001110100111;
		16'b1000011011010011: color_data = 12'b001110100111;
		16'b1000011011010100: color_data = 12'b001110100111;
		16'b1000011011010101: color_data = 12'b001110100111;
		16'b1000011011010110: color_data = 12'b001110100111;
		16'b1000011011110110: color_data = 12'b001110100111;
		16'b1000011011110111: color_data = 12'b001110100111;
		16'b1000011011111000: color_data = 12'b001110100111;
		16'b1000011011111001: color_data = 12'b001110100111;
		16'b1000011011111010: color_data = 12'b001110100111;
		16'b1000011011111011: color_data = 12'b001110100111;
		16'b1000011011111100: color_data = 12'b001110100111;
		16'b1000011011111101: color_data = 12'b001110100111;
		16'b1000011011111110: color_data = 12'b001110100111;
		16'b1000011011111111: color_data = 12'b001110100111;
		16'b1000011100000000: color_data = 12'b001110100111;
		16'b1000011100000001: color_data = 12'b001110100111;
		16'b1000011100011010: color_data = 12'b001110100111;
		16'b1000011100011011: color_data = 12'b001110100111;
		16'b1000011100011100: color_data = 12'b001110100111;
		16'b1000011100011101: color_data = 12'b001110100111;
		16'b1000011100011110: color_data = 12'b001110100111;
		16'b1000011100011111: color_data = 12'b001110100111;
		16'b1000011100100000: color_data = 12'b001110100111;
		16'b1000011100100001: color_data = 12'b001110100111;
		16'b1000011100100010: color_data = 12'b001110100111;
		16'b1000011100100011: color_data = 12'b001110100111;
		16'b1000011100100100: color_data = 12'b001110100111;
		16'b1000011100100101: color_data = 12'b001110100111;
		16'b1000011100100110: color_data = 12'b001110100111;
		16'b1000011100101101: color_data = 12'b001110100111;
		16'b1000011100101110: color_data = 12'b001110100111;
		16'b1000011100101111: color_data = 12'b001110100111;
		16'b1000011100110000: color_data = 12'b001110100111;
		16'b1000011100110001: color_data = 12'b001110100111;
		16'b1000011100110010: color_data = 12'b001110100111;
		16'b1000011100110011: color_data = 12'b001110100111;
		16'b1000011100110100: color_data = 12'b001110100111;
		16'b1000011100110101: color_data = 12'b001110100111;
		16'b1000011100110110: color_data = 12'b001110100111;
		16'b1000011100110111: color_data = 12'b001110100111;
		16'b1000011100111000: color_data = 12'b001110100111;
		16'b1000011101000101: color_data = 12'b001110100111;
		16'b1000011101000110: color_data = 12'b001110100111;
		16'b1000011101000111: color_data = 12'b001110100111;
		16'b1000011101001000: color_data = 12'b001110100111;
		16'b1000011101001001: color_data = 12'b001110100111;
		16'b1000011101001010: color_data = 12'b001110100111;
		16'b1000011101001011: color_data = 12'b001110100111;
		16'b1000011101001100: color_data = 12'b001110100111;
		16'b1000011101001101: color_data = 12'b001110100111;
		16'b1000011101001110: color_data = 12'b001110100111;
		16'b1000011101001111: color_data = 12'b001110100111;
		16'b1000011101010000: color_data = 12'b001110100111;
		16'b1000011101010001: color_data = 12'b001110100111;
		16'b1000011101011000: color_data = 12'b001110100111;
		16'b1000011101011001: color_data = 12'b001110100111;
		16'b1000011101011010: color_data = 12'b001110100111;
		16'b1000011101011011: color_data = 12'b001110100111;
		16'b1000011101011100: color_data = 12'b001110100111;
		16'b1000011101011101: color_data = 12'b001110100111;
		16'b1000011101011110: color_data = 12'b001110100111;
		16'b1000011101011111: color_data = 12'b001110100111;
		16'b1000011101100000: color_data = 12'b001110100111;
		16'b1000011101100001: color_data = 12'b001110100111;
		16'b1000011101100010: color_data = 12'b001110100111;
		16'b1000011101100011: color_data = 12'b001110100111;
		16'b1000011101110000: color_data = 12'b001110100111;
		16'b1000011101110001: color_data = 12'b001110100111;
		16'b1000011101110010: color_data = 12'b001110100111;
		16'b1000011101110011: color_data = 12'b001110100111;
		16'b1000011101110100: color_data = 12'b001110100111;
		16'b1000011101110101: color_data = 12'b001110100111;
		16'b1000011101110110: color_data = 12'b001110100111;
		16'b1000011101110111: color_data = 12'b001110100111;
		16'b1000011101111000: color_data = 12'b001110100111;
		16'b1000011101111001: color_data = 12'b001110100111;
		16'b1000011101111010: color_data = 12'b001110100111;
		16'b1000011101111011: color_data = 12'b001110100111;
		16'b1000100000000000: color_data = 12'b001110100111;
		16'b1000100000000001: color_data = 12'b001110100111;
		16'b1000100000000010: color_data = 12'b001110100111;
		16'b1000100000000011: color_data = 12'b001110100111;
		16'b1000100000000100: color_data = 12'b001110100111;
		16'b1000100000000101: color_data = 12'b001110100111;
		16'b1000100000000110: color_data = 12'b001110100111;
		16'b1000100000000111: color_data = 12'b001110100111;
		16'b1000100000001000: color_data = 12'b001110100111;
		16'b1000100000001001: color_data = 12'b001110100111;
		16'b1000100000001010: color_data = 12'b001110100111;
		16'b1000100000001011: color_data = 12'b001110100111;
		16'b1000100000001100: color_data = 12'b001110100111;
		16'b1000100000101011: color_data = 12'b001110100111;
		16'b1000100000101100: color_data = 12'b001110100111;
		16'b1000100000101101: color_data = 12'b001110100111;
		16'b1000100000101110: color_data = 12'b001110100111;
		16'b1000100000101111: color_data = 12'b001110100111;
		16'b1000100000110000: color_data = 12'b001110100111;
		16'b1000100000110001: color_data = 12'b001110100111;
		16'b1000100000110010: color_data = 12'b001110100111;
		16'b1000100000110011: color_data = 12'b001110100111;
		16'b1000100000110100: color_data = 12'b001110100111;
		16'b1000100000110101: color_data = 12'b001110100111;
		16'b1000100000110110: color_data = 12'b001110100111;
		16'b1000100000110111: color_data = 12'b001110100111;
		16'b1000100001000100: color_data = 12'b001110100111;
		16'b1000100001000101: color_data = 12'b001110100111;
		16'b1000100001000110: color_data = 12'b001110100111;
		16'b1000100001000111: color_data = 12'b001110100111;
		16'b1000100001001000: color_data = 12'b001110100111;
		16'b1000100001001001: color_data = 12'b001110100111;
		16'b1000100001001010: color_data = 12'b001110100111;
		16'b1000100001001011: color_data = 12'b001110100111;
		16'b1000100001001100: color_data = 12'b001110100111;
		16'b1000100001001101: color_data = 12'b001110100111;
		16'b1000100001001110: color_data = 12'b001110100111;
		16'b1000100001001111: color_data = 12'b001110100111;
		16'b1000100001011100: color_data = 12'b001110100111;
		16'b1000100001011101: color_data = 12'b001110100111;
		16'b1000100001011110: color_data = 12'b001110100111;
		16'b1000100001011111: color_data = 12'b001110100111;
		16'b1000100001100000: color_data = 12'b001110100111;
		16'b1000100001100001: color_data = 12'b001110100111;
		16'b1000100001100010: color_data = 12'b001110100111;
		16'b1000100001100011: color_data = 12'b001110100111;
		16'b1000100001100100: color_data = 12'b001110100111;
		16'b1000100001100101: color_data = 12'b001110100111;
		16'b1000100001100110: color_data = 12'b001110100111;
		16'b1000100001100111: color_data = 12'b001110100111;
		16'b1000100001101000: color_data = 12'b001110100111;
		16'b1000100001110101: color_data = 12'b001110100111;
		16'b1000100001110110: color_data = 12'b001110100111;
		16'b1000100001110111: color_data = 12'b001110100111;
		16'b1000100001111000: color_data = 12'b001110100111;
		16'b1000100001111001: color_data = 12'b001110100111;
		16'b1000100001111010: color_data = 12'b001110100111;
		16'b1000100001111011: color_data = 12'b001110100111;
		16'b1000100001111100: color_data = 12'b001110100111;
		16'b1000100001111101: color_data = 12'b001110100111;
		16'b1000100001111110: color_data = 12'b001110100111;
		16'b1000100001111111: color_data = 12'b001110100111;
		16'b1000100010000000: color_data = 12'b001110100111;
		16'b1000100010001101: color_data = 12'b001110100111;
		16'b1000100010001110: color_data = 12'b001110100111;
		16'b1000100010001111: color_data = 12'b001110100111;
		16'b1000100010010000: color_data = 12'b001110100111;
		16'b1000100010010001: color_data = 12'b001110100111;
		16'b1000100010010010: color_data = 12'b001110100111;
		16'b1000100010010011: color_data = 12'b001110100111;
		16'b1000100010010100: color_data = 12'b001110100111;
		16'b1000100010010101: color_data = 12'b001110100111;
		16'b1000100010010110: color_data = 12'b001110100111;
		16'b1000100010010111: color_data = 12'b001110100111;
		16'b1000100010011000: color_data = 12'b001110100111;
		16'b1000100010011001: color_data = 12'b001110100111;
		16'b1000100010100000: color_data = 12'b001110100111;
		16'b1000100010100001: color_data = 12'b001110100111;
		16'b1000100010100010: color_data = 12'b001110100111;
		16'b1000100010100011: color_data = 12'b001110100111;
		16'b1000100010100100: color_data = 12'b001110100111;
		16'b1000100010100101: color_data = 12'b001110100111;
		16'b1000100010100110: color_data = 12'b001110100111;
		16'b1000100010100111: color_data = 12'b001110100111;
		16'b1000100010101000: color_data = 12'b001110100111;
		16'b1000100010101001: color_data = 12'b001110100111;
		16'b1000100010101010: color_data = 12'b001110100111;
		16'b1000100010101011: color_data = 12'b001110100111;
		16'b1000100010111000: color_data = 12'b001110100111;
		16'b1000100010111001: color_data = 12'b001110100111;
		16'b1000100010111010: color_data = 12'b001110100111;
		16'b1000100010111011: color_data = 12'b001110100111;
		16'b1000100010111100: color_data = 12'b001110100111;
		16'b1000100010111101: color_data = 12'b001110100111;
		16'b1000100010111110: color_data = 12'b001110100111;
		16'b1000100010111111: color_data = 12'b001110100111;
		16'b1000100011000000: color_data = 12'b001110100111;
		16'b1000100011000001: color_data = 12'b001110100111;
		16'b1000100011000010: color_data = 12'b001110100111;
		16'b1000100011000011: color_data = 12'b001110100111;
		16'b1000100011000100: color_data = 12'b001110100111;
		16'b1000100011001011: color_data = 12'b001110100111;
		16'b1000100011001100: color_data = 12'b001110100111;
		16'b1000100011001101: color_data = 12'b001110100111;
		16'b1000100011001110: color_data = 12'b001110100111;
		16'b1000100011001111: color_data = 12'b001110100111;
		16'b1000100011010000: color_data = 12'b001110100111;
		16'b1000100011010001: color_data = 12'b001110100111;
		16'b1000100011010010: color_data = 12'b001110100111;
		16'b1000100011010011: color_data = 12'b001110100111;
		16'b1000100011010100: color_data = 12'b001110100111;
		16'b1000100011010101: color_data = 12'b001110100111;
		16'b1000100011010110: color_data = 12'b001110100111;
		16'b1000100011110110: color_data = 12'b001110100111;
		16'b1000100011110111: color_data = 12'b001110100111;
		16'b1000100011111000: color_data = 12'b001110100111;
		16'b1000100011111001: color_data = 12'b001110100111;
		16'b1000100011111010: color_data = 12'b001110100111;
		16'b1000100011111011: color_data = 12'b001110100111;
		16'b1000100011111100: color_data = 12'b001110100111;
		16'b1000100011111101: color_data = 12'b001110100111;
		16'b1000100011111110: color_data = 12'b001110100111;
		16'b1000100011111111: color_data = 12'b001110100111;
		16'b1000100100000000: color_data = 12'b001110100111;
		16'b1000100100000001: color_data = 12'b001110100111;
		16'b1000100100011010: color_data = 12'b001110100111;
		16'b1000100100011011: color_data = 12'b001110100111;
		16'b1000100100011100: color_data = 12'b001110100111;
		16'b1000100100011101: color_data = 12'b001110100111;
		16'b1000100100011110: color_data = 12'b001110100111;
		16'b1000100100011111: color_data = 12'b001110100111;
		16'b1000100100100000: color_data = 12'b001110100111;
		16'b1000100100100001: color_data = 12'b001110100111;
		16'b1000100100100010: color_data = 12'b001110100111;
		16'b1000100100100011: color_data = 12'b001110100111;
		16'b1000100100100100: color_data = 12'b001110100111;
		16'b1000100100100101: color_data = 12'b001110100111;
		16'b1000100100100110: color_data = 12'b001110100111;
		16'b1000100100101101: color_data = 12'b001110100111;
		16'b1000100100101110: color_data = 12'b001110100111;
		16'b1000100100101111: color_data = 12'b001110100111;
		16'b1000100100110000: color_data = 12'b001110100111;
		16'b1000100100110001: color_data = 12'b001110100111;
		16'b1000100100110010: color_data = 12'b001110100111;
		16'b1000100100110011: color_data = 12'b001110100111;
		16'b1000100100110100: color_data = 12'b001110100111;
		16'b1000100100110101: color_data = 12'b001110100111;
		16'b1000100100110110: color_data = 12'b001110100111;
		16'b1000100100110111: color_data = 12'b001110100111;
		16'b1000100100111000: color_data = 12'b001110100111;
		16'b1000100101000101: color_data = 12'b001110100111;
		16'b1000100101000110: color_data = 12'b001110100111;
		16'b1000100101000111: color_data = 12'b001110100111;
		16'b1000100101001000: color_data = 12'b001110100111;
		16'b1000100101001001: color_data = 12'b001110100111;
		16'b1000100101001010: color_data = 12'b001110100111;
		16'b1000100101001011: color_data = 12'b001110100111;
		16'b1000100101001100: color_data = 12'b001110100111;
		16'b1000100101001101: color_data = 12'b001110100111;
		16'b1000100101001110: color_data = 12'b001110100111;
		16'b1000100101001111: color_data = 12'b001110100111;
		16'b1000100101010000: color_data = 12'b001110100111;
		16'b1000100101010001: color_data = 12'b001110100111;
		16'b1000100101011000: color_data = 12'b001110100111;
		16'b1000100101011001: color_data = 12'b001110100111;
		16'b1000100101011010: color_data = 12'b001110100111;
		16'b1000100101011011: color_data = 12'b001110100111;
		16'b1000100101011100: color_data = 12'b001110100111;
		16'b1000100101011101: color_data = 12'b001110100111;
		16'b1000100101011110: color_data = 12'b001110100111;
		16'b1000100101011111: color_data = 12'b001110100111;
		16'b1000100101100000: color_data = 12'b001110100111;
		16'b1000100101100001: color_data = 12'b001110100111;
		16'b1000100101100010: color_data = 12'b001110100111;
		16'b1000100101100011: color_data = 12'b001110100111;
		16'b1000100101110000: color_data = 12'b001110100111;
		16'b1000100101110001: color_data = 12'b001110100111;
		16'b1000100101110010: color_data = 12'b001110100111;
		16'b1000100101110011: color_data = 12'b001110100111;
		16'b1000100101110100: color_data = 12'b001110100111;
		16'b1000100101110101: color_data = 12'b001110100111;
		16'b1000100101110110: color_data = 12'b001110100111;
		16'b1000100101110111: color_data = 12'b001110100111;
		16'b1000100101111000: color_data = 12'b001110100111;
		16'b1000100101111001: color_data = 12'b001110100111;
		16'b1000100101111010: color_data = 12'b001110100111;
		16'b1000100101111011: color_data = 12'b001110100111;
		16'b1000101000000000: color_data = 12'b001110100111;
		16'b1000101000000001: color_data = 12'b001110100111;
		16'b1000101000000010: color_data = 12'b001110100111;
		16'b1000101000000011: color_data = 12'b001110100111;
		16'b1000101000000100: color_data = 12'b001110100111;
		16'b1000101000000101: color_data = 12'b001110100111;
		16'b1000101000000110: color_data = 12'b001110100111;
		16'b1000101000000111: color_data = 12'b001110100111;
		16'b1000101000001000: color_data = 12'b001110100111;
		16'b1000101000001001: color_data = 12'b001110100111;
		16'b1000101000001010: color_data = 12'b001110100111;
		16'b1000101000001011: color_data = 12'b001110100111;
		16'b1000101000001100: color_data = 12'b001110100111;
		16'b1000101000101011: color_data = 12'b001110100111;
		16'b1000101000101100: color_data = 12'b001110100111;
		16'b1000101000101101: color_data = 12'b001110100111;
		16'b1000101000101110: color_data = 12'b001110100111;
		16'b1000101000101111: color_data = 12'b001110100111;
		16'b1000101000110000: color_data = 12'b001110100111;
		16'b1000101000110001: color_data = 12'b001110100111;
		16'b1000101000110010: color_data = 12'b001110100111;
		16'b1000101000110011: color_data = 12'b001110100111;
		16'b1000101000110100: color_data = 12'b001110100111;
		16'b1000101000110101: color_data = 12'b001110100111;
		16'b1000101000110110: color_data = 12'b001110100111;
		16'b1000101000110111: color_data = 12'b001110100111;
		16'b1000101001000100: color_data = 12'b001110100111;
		16'b1000101001000101: color_data = 12'b001110100111;
		16'b1000101001000110: color_data = 12'b001110100111;
		16'b1000101001000111: color_data = 12'b001110100111;
		16'b1000101001001000: color_data = 12'b001110100111;
		16'b1000101001001001: color_data = 12'b001110100111;
		16'b1000101001001010: color_data = 12'b001110100111;
		16'b1000101001001011: color_data = 12'b001110100111;
		16'b1000101001001100: color_data = 12'b001110100111;
		16'b1000101001001101: color_data = 12'b001110100111;
		16'b1000101001001110: color_data = 12'b001110100111;
		16'b1000101001001111: color_data = 12'b001110100111;
		16'b1000101001011100: color_data = 12'b001110100111;
		16'b1000101001011101: color_data = 12'b001110100111;
		16'b1000101001011110: color_data = 12'b001110100111;
		16'b1000101001011111: color_data = 12'b001110100111;
		16'b1000101001100000: color_data = 12'b001110100111;
		16'b1000101001100001: color_data = 12'b001110100111;
		16'b1000101001100010: color_data = 12'b001110100111;
		16'b1000101001100011: color_data = 12'b001110100111;
		16'b1000101001100100: color_data = 12'b001110100111;
		16'b1000101001100101: color_data = 12'b001110100111;
		16'b1000101001100110: color_data = 12'b001110100111;
		16'b1000101001100111: color_data = 12'b001110100111;
		16'b1000101001101000: color_data = 12'b001110100111;
		16'b1000101001110101: color_data = 12'b001110100111;
		16'b1000101001110110: color_data = 12'b001110100111;
		16'b1000101001110111: color_data = 12'b001110100111;
		16'b1000101001111000: color_data = 12'b001110100111;
		16'b1000101001111001: color_data = 12'b001110100111;
		16'b1000101001111010: color_data = 12'b001110100111;
		16'b1000101001111011: color_data = 12'b001110100111;
		16'b1000101001111100: color_data = 12'b001110100111;
		16'b1000101001111101: color_data = 12'b001110100111;
		16'b1000101001111110: color_data = 12'b001110100111;
		16'b1000101001111111: color_data = 12'b001110100111;
		16'b1000101010000000: color_data = 12'b001110100111;
		16'b1000101010001101: color_data = 12'b001110100111;
		16'b1000101010001110: color_data = 12'b001110100111;
		16'b1000101010001111: color_data = 12'b001110100111;
		16'b1000101010010000: color_data = 12'b001110100111;
		16'b1000101010010001: color_data = 12'b001110100111;
		16'b1000101010010010: color_data = 12'b001110100111;
		16'b1000101010010011: color_data = 12'b001110100111;
		16'b1000101010010100: color_data = 12'b001110100111;
		16'b1000101010010101: color_data = 12'b001110100111;
		16'b1000101010010110: color_data = 12'b001110100111;
		16'b1000101010010111: color_data = 12'b001110100111;
		16'b1000101010011000: color_data = 12'b001110100111;
		16'b1000101010011001: color_data = 12'b001110100111;
		16'b1000101010100000: color_data = 12'b001110100111;
		16'b1000101010100001: color_data = 12'b001110100111;
		16'b1000101010100010: color_data = 12'b001110100111;
		16'b1000101010100011: color_data = 12'b001110100111;
		16'b1000101010100100: color_data = 12'b001110100111;
		16'b1000101010100101: color_data = 12'b001110100111;
		16'b1000101010100110: color_data = 12'b001110100111;
		16'b1000101010100111: color_data = 12'b001110100111;
		16'b1000101010101000: color_data = 12'b001110100111;
		16'b1000101010101001: color_data = 12'b001110100111;
		16'b1000101010101010: color_data = 12'b001110100111;
		16'b1000101010101011: color_data = 12'b001110100111;
		16'b1000101010111000: color_data = 12'b001110100111;
		16'b1000101010111001: color_data = 12'b001110100111;
		16'b1000101010111010: color_data = 12'b001110100111;
		16'b1000101010111011: color_data = 12'b001110100111;
		16'b1000101010111100: color_data = 12'b001110100111;
		16'b1000101010111101: color_data = 12'b001110100111;
		16'b1000101010111110: color_data = 12'b001110100111;
		16'b1000101010111111: color_data = 12'b001110100111;
		16'b1000101011000000: color_data = 12'b001110100111;
		16'b1000101011000001: color_data = 12'b001110100111;
		16'b1000101011000010: color_data = 12'b001110100111;
		16'b1000101011000011: color_data = 12'b001110100111;
		16'b1000101011000100: color_data = 12'b001110100111;
		16'b1000101011001011: color_data = 12'b001110100111;
		16'b1000101011001100: color_data = 12'b001110100111;
		16'b1000101011001101: color_data = 12'b001110100111;
		16'b1000101011001110: color_data = 12'b001110100111;
		16'b1000101011001111: color_data = 12'b001110100111;
		16'b1000101011010000: color_data = 12'b001110100111;
		16'b1000101011010001: color_data = 12'b001110100111;
		16'b1000101011010010: color_data = 12'b001110100111;
		16'b1000101011010011: color_data = 12'b001110100111;
		16'b1000101011010100: color_data = 12'b001110100111;
		16'b1000101011010101: color_data = 12'b001110100111;
		16'b1000101011010110: color_data = 12'b001110100111;
		16'b1000101011110110: color_data = 12'b001110100111;
		16'b1000101011110111: color_data = 12'b001110100111;
		16'b1000101011111000: color_data = 12'b001110100111;
		16'b1000101011111001: color_data = 12'b001110100111;
		16'b1000101011111010: color_data = 12'b001110100111;
		16'b1000101011111011: color_data = 12'b001110100111;
		16'b1000101011111100: color_data = 12'b001110100111;
		16'b1000101011111101: color_data = 12'b001110100111;
		16'b1000101011111110: color_data = 12'b001110100111;
		16'b1000101011111111: color_data = 12'b001110100111;
		16'b1000101100000000: color_data = 12'b001110100111;
		16'b1000101100000001: color_data = 12'b001110100111;
		16'b1000101100011010: color_data = 12'b001110100111;
		16'b1000101100011011: color_data = 12'b001110100111;
		16'b1000101100011100: color_data = 12'b001110100111;
		16'b1000101100011101: color_data = 12'b001110100111;
		16'b1000101100011110: color_data = 12'b001110100111;
		16'b1000101100011111: color_data = 12'b001110100111;
		16'b1000101100100000: color_data = 12'b001110100111;
		16'b1000101100100001: color_data = 12'b001110100111;
		16'b1000101100100010: color_data = 12'b001110100111;
		16'b1000101100100011: color_data = 12'b001110100111;
		16'b1000101100100100: color_data = 12'b001110100111;
		16'b1000101100100101: color_data = 12'b001110100111;
		16'b1000101100100110: color_data = 12'b001110100111;
		16'b1000101100101101: color_data = 12'b001110100111;
		16'b1000101100101110: color_data = 12'b001110100111;
		16'b1000101100101111: color_data = 12'b001110100111;
		16'b1000101100110000: color_data = 12'b001110100111;
		16'b1000101100110001: color_data = 12'b001110100111;
		16'b1000101100110010: color_data = 12'b001110100111;
		16'b1000101100110011: color_data = 12'b001110100111;
		16'b1000101100110100: color_data = 12'b001110100111;
		16'b1000101100110101: color_data = 12'b001110100111;
		16'b1000101100110110: color_data = 12'b001110100111;
		16'b1000101100110111: color_data = 12'b001110100111;
		16'b1000101100111000: color_data = 12'b001110100111;
		16'b1000101101000101: color_data = 12'b001110100111;
		16'b1000101101000110: color_data = 12'b001110100111;
		16'b1000101101000111: color_data = 12'b001110100111;
		16'b1000101101001000: color_data = 12'b001110100111;
		16'b1000101101001001: color_data = 12'b001110100111;
		16'b1000101101001010: color_data = 12'b001110100111;
		16'b1000101101001011: color_data = 12'b001110100111;
		16'b1000101101001100: color_data = 12'b001110100111;
		16'b1000101101001101: color_data = 12'b001110100111;
		16'b1000101101001110: color_data = 12'b001110100111;
		16'b1000101101001111: color_data = 12'b001110100111;
		16'b1000101101010000: color_data = 12'b001110100111;
		16'b1000101101010001: color_data = 12'b001110100111;
		16'b1000101101011000: color_data = 12'b001110100111;
		16'b1000101101011001: color_data = 12'b001110100111;
		16'b1000101101011010: color_data = 12'b001110100111;
		16'b1000101101011011: color_data = 12'b001110100111;
		16'b1000101101011100: color_data = 12'b001110100111;
		16'b1000101101011101: color_data = 12'b001110100111;
		16'b1000101101011110: color_data = 12'b001110100111;
		16'b1000101101011111: color_data = 12'b001110100111;
		16'b1000101101100000: color_data = 12'b001110100111;
		16'b1000101101100001: color_data = 12'b001110100111;
		16'b1000101101100010: color_data = 12'b001110100111;
		16'b1000101101100011: color_data = 12'b001110100111;
		16'b1000101101110000: color_data = 12'b001110100111;
		16'b1000101101110001: color_data = 12'b001110100111;
		16'b1000101101110010: color_data = 12'b001110100111;
		16'b1000101101110011: color_data = 12'b001110100111;
		16'b1000101101110100: color_data = 12'b001110100111;
		16'b1000101101110101: color_data = 12'b001110100111;
		16'b1000101101110110: color_data = 12'b001110100111;
		16'b1000101101110111: color_data = 12'b001110100111;
		16'b1000101101111000: color_data = 12'b001110100111;
		16'b1000101101111001: color_data = 12'b001110100111;
		16'b1000101101111010: color_data = 12'b001110100111;
		16'b1000101101111011: color_data = 12'b001110100111;
		16'b1000110000000000: color_data = 12'b001110100111;
		16'b1000110000000001: color_data = 12'b001110100111;
		16'b1000110000000010: color_data = 12'b001110100111;
		16'b1000110000000011: color_data = 12'b001110100111;
		16'b1000110000000100: color_data = 12'b001110100111;
		16'b1000110000000101: color_data = 12'b001110100111;
		16'b1000110000000110: color_data = 12'b001110100111;
		16'b1000110000000111: color_data = 12'b001110100111;
		16'b1000110000001000: color_data = 12'b001110100111;
		16'b1000110000001001: color_data = 12'b001110100111;
		16'b1000110000001010: color_data = 12'b001110100111;
		16'b1000110000001011: color_data = 12'b001110100111;
		16'b1000110000001100: color_data = 12'b001110100111;
		16'b1000110000101011: color_data = 12'b001110100111;
		16'b1000110000101100: color_data = 12'b001110100111;
		16'b1000110000101101: color_data = 12'b001110100111;
		16'b1000110000101110: color_data = 12'b001110100111;
		16'b1000110000101111: color_data = 12'b001110100111;
		16'b1000110000110000: color_data = 12'b001110100111;
		16'b1000110000110001: color_data = 12'b001110100111;
		16'b1000110000110010: color_data = 12'b001110100111;
		16'b1000110000110011: color_data = 12'b001110100111;
		16'b1000110000110100: color_data = 12'b001110100111;
		16'b1000110000110101: color_data = 12'b001110100111;
		16'b1000110000110110: color_data = 12'b001110100111;
		16'b1000110000110111: color_data = 12'b001110100111;
		16'b1000110001000100: color_data = 12'b001110100111;
		16'b1000110001000101: color_data = 12'b001110100111;
		16'b1000110001000110: color_data = 12'b001110100111;
		16'b1000110001000111: color_data = 12'b001110100111;
		16'b1000110001001000: color_data = 12'b001110100111;
		16'b1000110001001001: color_data = 12'b001110100111;
		16'b1000110001001010: color_data = 12'b001110100111;
		16'b1000110001001011: color_data = 12'b001110100111;
		16'b1000110001001100: color_data = 12'b001110100111;
		16'b1000110001001101: color_data = 12'b001110100111;
		16'b1000110001001110: color_data = 12'b001110100111;
		16'b1000110001001111: color_data = 12'b001110100111;
		16'b1000110001011100: color_data = 12'b001110100111;
		16'b1000110001011101: color_data = 12'b001110100111;
		16'b1000110001011110: color_data = 12'b001110100111;
		16'b1000110001011111: color_data = 12'b001110100111;
		16'b1000110001100000: color_data = 12'b001110100111;
		16'b1000110001100001: color_data = 12'b001110100111;
		16'b1000110001100010: color_data = 12'b001110100111;
		16'b1000110001100011: color_data = 12'b001110100111;
		16'b1000110001100100: color_data = 12'b001110100111;
		16'b1000110001100101: color_data = 12'b001110100111;
		16'b1000110001100110: color_data = 12'b001110100111;
		16'b1000110001100111: color_data = 12'b001110100111;
		16'b1000110001101000: color_data = 12'b001110100111;
		16'b1000110001110101: color_data = 12'b001110100111;
		16'b1000110001110110: color_data = 12'b001110100111;
		16'b1000110001110111: color_data = 12'b001110100111;
		16'b1000110001111000: color_data = 12'b001110100111;
		16'b1000110001111001: color_data = 12'b001110100111;
		16'b1000110001111010: color_data = 12'b001110100111;
		16'b1000110001111011: color_data = 12'b001110100111;
		16'b1000110001111100: color_data = 12'b001110100111;
		16'b1000110001111101: color_data = 12'b001110100111;
		16'b1000110001111110: color_data = 12'b001110100111;
		16'b1000110001111111: color_data = 12'b001110100111;
		16'b1000110010000000: color_data = 12'b001110100111;
		16'b1000110010001101: color_data = 12'b001110100111;
		16'b1000110010001110: color_data = 12'b001110100111;
		16'b1000110010001111: color_data = 12'b001110100111;
		16'b1000110010010000: color_data = 12'b001110100111;
		16'b1000110010010001: color_data = 12'b001110100111;
		16'b1000110010010010: color_data = 12'b001110100111;
		16'b1000110010010011: color_data = 12'b001110100111;
		16'b1000110010010100: color_data = 12'b001110100111;
		16'b1000110010010101: color_data = 12'b001110100111;
		16'b1000110010010110: color_data = 12'b001110100111;
		16'b1000110010010111: color_data = 12'b001110100111;
		16'b1000110010011000: color_data = 12'b001110100111;
		16'b1000110010011001: color_data = 12'b001110100111;
		16'b1000110010100000: color_data = 12'b001110100111;
		16'b1000110010100001: color_data = 12'b001110100111;
		16'b1000110010100010: color_data = 12'b001110100111;
		16'b1000110010100011: color_data = 12'b001110100111;
		16'b1000110010100100: color_data = 12'b001110100111;
		16'b1000110010100101: color_data = 12'b001110100111;
		16'b1000110010100110: color_data = 12'b001110100111;
		16'b1000110010100111: color_data = 12'b001110100111;
		16'b1000110010101000: color_data = 12'b001110100111;
		16'b1000110010101001: color_data = 12'b001110100111;
		16'b1000110010101010: color_data = 12'b001110100111;
		16'b1000110010101011: color_data = 12'b001110100111;
		16'b1000110010111000: color_data = 12'b001110100111;
		16'b1000110010111001: color_data = 12'b001110100111;
		16'b1000110010111010: color_data = 12'b001110100111;
		16'b1000110010111011: color_data = 12'b001110100111;
		16'b1000110010111100: color_data = 12'b001110100111;
		16'b1000110010111101: color_data = 12'b001110100111;
		16'b1000110010111110: color_data = 12'b001110100111;
		16'b1000110010111111: color_data = 12'b001110100111;
		16'b1000110011000000: color_data = 12'b001110100111;
		16'b1000110011000001: color_data = 12'b001110100111;
		16'b1000110011000010: color_data = 12'b001110100111;
		16'b1000110011000011: color_data = 12'b001110100111;
		16'b1000110011000100: color_data = 12'b001110100111;
		16'b1000110011001011: color_data = 12'b001110100111;
		16'b1000110011001100: color_data = 12'b001110100111;
		16'b1000110011001101: color_data = 12'b001110100111;
		16'b1000110011001110: color_data = 12'b001110100111;
		16'b1000110011001111: color_data = 12'b001110100111;
		16'b1000110011010000: color_data = 12'b001110100111;
		16'b1000110011010001: color_data = 12'b001110100111;
		16'b1000110011010010: color_data = 12'b001110100111;
		16'b1000110011010011: color_data = 12'b001110100111;
		16'b1000110011010100: color_data = 12'b001110100111;
		16'b1000110011010101: color_data = 12'b001110100111;
		16'b1000110011010110: color_data = 12'b001110100111;
		16'b1000110011110110: color_data = 12'b001110100111;
		16'b1000110011110111: color_data = 12'b001110100111;
		16'b1000110011111000: color_data = 12'b001110100111;
		16'b1000110011111001: color_data = 12'b001110100111;
		16'b1000110011111010: color_data = 12'b001110100111;
		16'b1000110011111011: color_data = 12'b001110100111;
		16'b1000110011111100: color_data = 12'b001110100111;
		16'b1000110011111101: color_data = 12'b001110100111;
		16'b1000110011111110: color_data = 12'b001110100111;
		16'b1000110011111111: color_data = 12'b001110100111;
		16'b1000110100000000: color_data = 12'b001110100111;
		16'b1000110100000001: color_data = 12'b001110100111;
		16'b1000110100011010: color_data = 12'b001110100111;
		16'b1000110100011011: color_data = 12'b001110100111;
		16'b1000110100011100: color_data = 12'b001110100111;
		16'b1000110100011101: color_data = 12'b001110100111;
		16'b1000110100011110: color_data = 12'b001110100111;
		16'b1000110100011111: color_data = 12'b001110100111;
		16'b1000110100100000: color_data = 12'b001110100111;
		16'b1000110100100001: color_data = 12'b001110100111;
		16'b1000110100100010: color_data = 12'b001110100111;
		16'b1000110100100011: color_data = 12'b001110100111;
		16'b1000110100100100: color_data = 12'b001110100111;
		16'b1000110100100101: color_data = 12'b001110100111;
		16'b1000110100100110: color_data = 12'b001110100111;
		16'b1000110100101101: color_data = 12'b001110100111;
		16'b1000110100101110: color_data = 12'b001110100111;
		16'b1000110100101111: color_data = 12'b001110100111;
		16'b1000110100110000: color_data = 12'b001110100111;
		16'b1000110100110001: color_data = 12'b001110100111;
		16'b1000110100110010: color_data = 12'b001110100111;
		16'b1000110100110011: color_data = 12'b001110100111;
		16'b1000110100110100: color_data = 12'b001110100111;
		16'b1000110100110101: color_data = 12'b001110100111;
		16'b1000110100110110: color_data = 12'b001110100111;
		16'b1000110100110111: color_data = 12'b001110100111;
		16'b1000110100111000: color_data = 12'b001110100111;
		16'b1000110101000101: color_data = 12'b001110100111;
		16'b1000110101000110: color_data = 12'b001110100111;
		16'b1000110101000111: color_data = 12'b001110100111;
		16'b1000110101001000: color_data = 12'b001110100111;
		16'b1000110101001001: color_data = 12'b001110100111;
		16'b1000110101001010: color_data = 12'b001110100111;
		16'b1000110101001011: color_data = 12'b001110100111;
		16'b1000110101001100: color_data = 12'b001110100111;
		16'b1000110101001101: color_data = 12'b001110100111;
		16'b1000110101001110: color_data = 12'b001110100111;
		16'b1000110101001111: color_data = 12'b001110100111;
		16'b1000110101010000: color_data = 12'b001110100111;
		16'b1000110101010001: color_data = 12'b001110100111;
		16'b1000110101011000: color_data = 12'b001110100111;
		16'b1000110101011001: color_data = 12'b001110100111;
		16'b1000110101011010: color_data = 12'b001110100111;
		16'b1000110101011011: color_data = 12'b001110100111;
		16'b1000110101011100: color_data = 12'b001110100111;
		16'b1000110101011101: color_data = 12'b001110100111;
		16'b1000110101011110: color_data = 12'b001110100111;
		16'b1000110101011111: color_data = 12'b001110100111;
		16'b1000110101100000: color_data = 12'b001110100111;
		16'b1000110101100001: color_data = 12'b001110100111;
		16'b1000110101100010: color_data = 12'b001110100111;
		16'b1000110101100011: color_data = 12'b001110100111;
		16'b1000110101110000: color_data = 12'b001110100111;
		16'b1000110101110001: color_data = 12'b001110100111;
		16'b1000110101110010: color_data = 12'b001110100111;
		16'b1000110101110011: color_data = 12'b001110100111;
		16'b1000110101110100: color_data = 12'b001110100111;
		16'b1000110101110101: color_data = 12'b001110100111;
		16'b1000110101110110: color_data = 12'b001110100111;
		16'b1000110101110111: color_data = 12'b001110100111;
		16'b1000110101111000: color_data = 12'b001110100111;
		16'b1000110101111001: color_data = 12'b001110100111;
		16'b1000110101111010: color_data = 12'b001110100111;
		16'b1000110101111011: color_data = 12'b001110100111;
		16'b1000111000000000: color_data = 12'b001110100111;
		16'b1000111000000001: color_data = 12'b001110100111;
		16'b1000111000000010: color_data = 12'b001110100111;
		16'b1000111000000011: color_data = 12'b001110100111;
		16'b1000111000000100: color_data = 12'b001110100111;
		16'b1000111000000101: color_data = 12'b001110100111;
		16'b1000111000000110: color_data = 12'b001110100111;
		16'b1000111000000111: color_data = 12'b001110100111;
		16'b1000111000001000: color_data = 12'b001110100111;
		16'b1000111000001001: color_data = 12'b001110100111;
		16'b1000111000001010: color_data = 12'b001110100111;
		16'b1000111000001011: color_data = 12'b001110100111;
		16'b1000111000001100: color_data = 12'b001110100111;
		16'b1000111000101011: color_data = 12'b001110100111;
		16'b1000111000101100: color_data = 12'b001110100111;
		16'b1000111000101101: color_data = 12'b001110100111;
		16'b1000111000101110: color_data = 12'b001110100111;
		16'b1000111000101111: color_data = 12'b001110100111;
		16'b1000111000110000: color_data = 12'b001110100111;
		16'b1000111000110001: color_data = 12'b001110100111;
		16'b1000111000110010: color_data = 12'b001110100111;
		16'b1000111000110011: color_data = 12'b001110100111;
		16'b1000111000110100: color_data = 12'b001110100111;
		16'b1000111000110101: color_data = 12'b001110100111;
		16'b1000111000110110: color_data = 12'b001110100111;
		16'b1000111000110111: color_data = 12'b001110100111;
		16'b1000111001000100: color_data = 12'b001110100111;
		16'b1000111001000101: color_data = 12'b001110100111;
		16'b1000111001000110: color_data = 12'b001110100111;
		16'b1000111001000111: color_data = 12'b001110100111;
		16'b1000111001001000: color_data = 12'b001110100111;
		16'b1000111001001001: color_data = 12'b001110100111;
		16'b1000111001001010: color_data = 12'b001110100111;
		16'b1000111001001011: color_data = 12'b001110100111;
		16'b1000111001001100: color_data = 12'b001110100111;
		16'b1000111001001101: color_data = 12'b001110100111;
		16'b1000111001001110: color_data = 12'b001110100111;
		16'b1000111001001111: color_data = 12'b001110100111;
		16'b1000111001011100: color_data = 12'b001110100111;
		16'b1000111001011101: color_data = 12'b001110100111;
		16'b1000111001011110: color_data = 12'b001110100111;
		16'b1000111001011111: color_data = 12'b001110100111;
		16'b1000111001100000: color_data = 12'b001110100111;
		16'b1000111001100001: color_data = 12'b001110100111;
		16'b1000111001100010: color_data = 12'b001110100111;
		16'b1000111001100011: color_data = 12'b001110100111;
		16'b1000111001100100: color_data = 12'b001110100111;
		16'b1000111001100101: color_data = 12'b001110100111;
		16'b1000111001100110: color_data = 12'b001110100111;
		16'b1000111001100111: color_data = 12'b001110100111;
		16'b1000111001101000: color_data = 12'b001110100111;
		16'b1000111001110101: color_data = 12'b001110100111;
		16'b1000111001110110: color_data = 12'b001110100111;
		16'b1000111001110111: color_data = 12'b001110100111;
		16'b1000111001111000: color_data = 12'b001110100111;
		16'b1000111001111001: color_data = 12'b001110100111;
		16'b1000111001111010: color_data = 12'b001110100111;
		16'b1000111001111011: color_data = 12'b001110100111;
		16'b1000111001111100: color_data = 12'b001110100111;
		16'b1000111001111101: color_data = 12'b001110100111;
		16'b1000111001111110: color_data = 12'b001110100111;
		16'b1000111001111111: color_data = 12'b001110100111;
		16'b1000111010000000: color_data = 12'b001110100111;
		16'b1000111010001101: color_data = 12'b001110100111;
		16'b1000111010001110: color_data = 12'b001110100111;
		16'b1000111010001111: color_data = 12'b001110100111;
		16'b1000111010010000: color_data = 12'b001110100111;
		16'b1000111010010001: color_data = 12'b001110100111;
		16'b1000111010010010: color_data = 12'b001110100111;
		16'b1000111010010011: color_data = 12'b001110100111;
		16'b1000111010010100: color_data = 12'b001110100111;
		16'b1000111010010101: color_data = 12'b001110100111;
		16'b1000111010010110: color_data = 12'b001110100111;
		16'b1000111010010111: color_data = 12'b001110100111;
		16'b1000111010011000: color_data = 12'b001110100111;
		16'b1000111010011001: color_data = 12'b001110100111;
		16'b1000111010100000: color_data = 12'b001110100111;
		16'b1000111010100001: color_data = 12'b001110100111;
		16'b1000111010100010: color_data = 12'b001110100111;
		16'b1000111010100011: color_data = 12'b001110100111;
		16'b1000111010100100: color_data = 12'b001110100111;
		16'b1000111010100101: color_data = 12'b001110100111;
		16'b1000111010100110: color_data = 12'b001110100111;
		16'b1000111010100111: color_data = 12'b001110100111;
		16'b1000111010101000: color_data = 12'b001110100111;
		16'b1000111010101001: color_data = 12'b001110100111;
		16'b1000111010101010: color_data = 12'b001110100111;
		16'b1000111010101011: color_data = 12'b001110100111;
		16'b1000111010111000: color_data = 12'b001110100111;
		16'b1000111010111001: color_data = 12'b001110100111;
		16'b1000111010111010: color_data = 12'b001110100111;
		16'b1000111010111011: color_data = 12'b001110100111;
		16'b1000111010111100: color_data = 12'b001110100111;
		16'b1000111010111101: color_data = 12'b001110100111;
		16'b1000111010111110: color_data = 12'b001110100111;
		16'b1000111010111111: color_data = 12'b001110100111;
		16'b1000111011000000: color_data = 12'b001110100111;
		16'b1000111011000001: color_data = 12'b001110100111;
		16'b1000111011000010: color_data = 12'b001110100111;
		16'b1000111011000011: color_data = 12'b001110100111;
		16'b1000111011000100: color_data = 12'b001110100111;
		16'b1000111011001011: color_data = 12'b001110100111;
		16'b1000111011001100: color_data = 12'b001110100111;
		16'b1000111011001101: color_data = 12'b001110100111;
		16'b1000111011001110: color_data = 12'b001110100111;
		16'b1000111011001111: color_data = 12'b001110100111;
		16'b1000111011010000: color_data = 12'b001110100111;
		16'b1000111011010001: color_data = 12'b001110100111;
		16'b1000111011010010: color_data = 12'b001110100111;
		16'b1000111011010011: color_data = 12'b001110100111;
		16'b1000111011010100: color_data = 12'b001110100111;
		16'b1000111011010101: color_data = 12'b001110100111;
		16'b1000111011010110: color_data = 12'b001110100111;
		16'b1000111011110110: color_data = 12'b001110100111;
		16'b1000111011110111: color_data = 12'b001110100111;
		16'b1000111011111000: color_data = 12'b001110100111;
		16'b1000111011111001: color_data = 12'b001110100111;
		16'b1000111011111010: color_data = 12'b001110100111;
		16'b1000111011111011: color_data = 12'b001110100111;
		16'b1000111011111100: color_data = 12'b001110100111;
		16'b1000111011111101: color_data = 12'b001110100111;
		16'b1000111011111110: color_data = 12'b001110100111;
		16'b1000111011111111: color_data = 12'b001110100111;
		16'b1000111100000000: color_data = 12'b001110100111;
		16'b1000111100000001: color_data = 12'b001110100111;
		16'b1000111100011010: color_data = 12'b001110100111;
		16'b1000111100011011: color_data = 12'b001110100111;
		16'b1000111100011100: color_data = 12'b001110100111;
		16'b1000111100011101: color_data = 12'b001110100111;
		16'b1000111100011110: color_data = 12'b001110100111;
		16'b1000111100011111: color_data = 12'b001110100111;
		16'b1000111100100000: color_data = 12'b001110100111;
		16'b1000111100100001: color_data = 12'b001110100111;
		16'b1000111100100010: color_data = 12'b001110100111;
		16'b1000111100100011: color_data = 12'b001110100111;
		16'b1000111100100100: color_data = 12'b001110100111;
		16'b1000111100100101: color_data = 12'b001110100111;
		16'b1000111100100110: color_data = 12'b001110100111;
		16'b1000111100101101: color_data = 12'b001110100111;
		16'b1000111100101110: color_data = 12'b001110100111;
		16'b1000111100101111: color_data = 12'b001110100111;
		16'b1000111100110000: color_data = 12'b001110100111;
		16'b1000111100110001: color_data = 12'b001110100111;
		16'b1000111100110010: color_data = 12'b001110100111;
		16'b1000111100110011: color_data = 12'b001110100111;
		16'b1000111100110100: color_data = 12'b001110100111;
		16'b1000111100110101: color_data = 12'b001110100111;
		16'b1000111100110110: color_data = 12'b001110100111;
		16'b1000111100110111: color_data = 12'b001110100111;
		16'b1000111100111000: color_data = 12'b001110100111;
		16'b1000111101000101: color_data = 12'b001110100111;
		16'b1000111101000110: color_data = 12'b001110100111;
		16'b1000111101000111: color_data = 12'b001110100111;
		16'b1000111101001000: color_data = 12'b001110100111;
		16'b1000111101001001: color_data = 12'b001110100111;
		16'b1000111101001010: color_data = 12'b001110100111;
		16'b1000111101001011: color_data = 12'b001110100111;
		16'b1000111101001100: color_data = 12'b001110100111;
		16'b1000111101001101: color_data = 12'b001110100111;
		16'b1000111101001110: color_data = 12'b001110100111;
		16'b1000111101001111: color_data = 12'b001110100111;
		16'b1000111101010000: color_data = 12'b001110100111;
		16'b1000111101010001: color_data = 12'b001110100111;
		16'b1000111101011000: color_data = 12'b001110100111;
		16'b1000111101011001: color_data = 12'b001110100111;
		16'b1000111101011010: color_data = 12'b001110100111;
		16'b1000111101011011: color_data = 12'b001110100111;
		16'b1000111101011100: color_data = 12'b001110100111;
		16'b1000111101011101: color_data = 12'b001110100111;
		16'b1000111101011110: color_data = 12'b001110100111;
		16'b1000111101011111: color_data = 12'b001110100111;
		16'b1000111101100000: color_data = 12'b001110100111;
		16'b1000111101100001: color_data = 12'b001110100111;
		16'b1000111101100010: color_data = 12'b001110100111;
		16'b1000111101100011: color_data = 12'b001110100111;
		16'b1000111101110000: color_data = 12'b001110100111;
		16'b1000111101110001: color_data = 12'b001110100111;
		16'b1000111101110010: color_data = 12'b001110100111;
		16'b1000111101110011: color_data = 12'b001110100111;
		16'b1000111101110100: color_data = 12'b001110100111;
		16'b1000111101110101: color_data = 12'b001110100111;
		16'b1000111101110110: color_data = 12'b001110100111;
		16'b1000111101110111: color_data = 12'b001110100111;
		16'b1000111101111000: color_data = 12'b001110100111;
		16'b1000111101111001: color_data = 12'b001110100111;
		16'b1000111101111010: color_data = 12'b001110100111;
		16'b1000111101111011: color_data = 12'b001110100111;
		16'b1001000000000000: color_data = 12'b001110100111;
		16'b1001000000000001: color_data = 12'b001110100111;
		16'b1001000000000010: color_data = 12'b001110100111;
		16'b1001000000000011: color_data = 12'b001110100111;
		16'b1001000000000100: color_data = 12'b001110100111;
		16'b1001000000000101: color_data = 12'b001110100111;
		16'b1001000000000110: color_data = 12'b001110100111;
		16'b1001000000000111: color_data = 12'b001110100111;
		16'b1001000000001000: color_data = 12'b001110100111;
		16'b1001000000001001: color_data = 12'b001110100111;
		16'b1001000000001010: color_data = 12'b001110100111;
		16'b1001000000001011: color_data = 12'b001110100111;
		16'b1001000000001100: color_data = 12'b001110100111;
		16'b1001000000101011: color_data = 12'b001110100111;
		16'b1001000000101100: color_data = 12'b001110100111;
		16'b1001000000101101: color_data = 12'b001110100111;
		16'b1001000000101110: color_data = 12'b001110100111;
		16'b1001000000101111: color_data = 12'b001110100111;
		16'b1001000000110000: color_data = 12'b001110100111;
		16'b1001000000110001: color_data = 12'b001110100111;
		16'b1001000000110010: color_data = 12'b001110100111;
		16'b1001000000110011: color_data = 12'b001110100111;
		16'b1001000000110100: color_data = 12'b001110100111;
		16'b1001000000110101: color_data = 12'b001110100111;
		16'b1001000000110110: color_data = 12'b001110100111;
		16'b1001000000110111: color_data = 12'b001110100111;
		16'b1001000001000100: color_data = 12'b001110100111;
		16'b1001000001000101: color_data = 12'b001110100111;
		16'b1001000001000110: color_data = 12'b001110100111;
		16'b1001000001000111: color_data = 12'b001110100111;
		16'b1001000001001000: color_data = 12'b001110100111;
		16'b1001000001001001: color_data = 12'b001110100111;
		16'b1001000001001010: color_data = 12'b001110100111;
		16'b1001000001001011: color_data = 12'b001110100111;
		16'b1001000001001100: color_data = 12'b001110100111;
		16'b1001000001001101: color_data = 12'b001110100111;
		16'b1001000001001110: color_data = 12'b001110100111;
		16'b1001000001001111: color_data = 12'b001110100111;
		16'b1001000001011100: color_data = 12'b001110100111;
		16'b1001000001011101: color_data = 12'b001110100111;
		16'b1001000001011110: color_data = 12'b001110100111;
		16'b1001000001011111: color_data = 12'b001110100111;
		16'b1001000001100000: color_data = 12'b001110100111;
		16'b1001000001100001: color_data = 12'b001110100111;
		16'b1001000001100010: color_data = 12'b001110100111;
		16'b1001000001100011: color_data = 12'b001110100111;
		16'b1001000001100100: color_data = 12'b001110100111;
		16'b1001000001100101: color_data = 12'b001110100111;
		16'b1001000001100110: color_data = 12'b001110100111;
		16'b1001000001100111: color_data = 12'b001110100111;
		16'b1001000001101000: color_data = 12'b001110100111;
		16'b1001000001110101: color_data = 12'b001110100111;
		16'b1001000001110110: color_data = 12'b001110100111;
		16'b1001000001110111: color_data = 12'b001110100111;
		16'b1001000001111000: color_data = 12'b001110100111;
		16'b1001000001111001: color_data = 12'b001110100111;
		16'b1001000001111010: color_data = 12'b001110100111;
		16'b1001000001111011: color_data = 12'b001110100111;
		16'b1001000001111100: color_data = 12'b001110100111;
		16'b1001000001111101: color_data = 12'b001110100111;
		16'b1001000001111110: color_data = 12'b001110100111;
		16'b1001000001111111: color_data = 12'b001110100111;
		16'b1001000010000000: color_data = 12'b001110100111;
		16'b1001000010001101: color_data = 12'b001110100111;
		16'b1001000010001110: color_data = 12'b001110100111;
		16'b1001000010001111: color_data = 12'b001110100111;
		16'b1001000010010000: color_data = 12'b001110100111;
		16'b1001000010010001: color_data = 12'b001110100111;
		16'b1001000010010010: color_data = 12'b001110100111;
		16'b1001000010010011: color_data = 12'b001110100111;
		16'b1001000010010100: color_data = 12'b001110100111;
		16'b1001000010010101: color_data = 12'b001110100111;
		16'b1001000010010110: color_data = 12'b001110100111;
		16'b1001000010010111: color_data = 12'b001110100111;
		16'b1001000010011000: color_data = 12'b001110100111;
		16'b1001000010011001: color_data = 12'b001110100111;
		16'b1001000010100000: color_data = 12'b001110100111;
		16'b1001000010100001: color_data = 12'b001110100111;
		16'b1001000010100010: color_data = 12'b001110100111;
		16'b1001000010100011: color_data = 12'b001110100111;
		16'b1001000010100100: color_data = 12'b001110100111;
		16'b1001000010100101: color_data = 12'b001110100111;
		16'b1001000010100110: color_data = 12'b001110100111;
		16'b1001000010100111: color_data = 12'b001110100111;
		16'b1001000010101000: color_data = 12'b001110100111;
		16'b1001000010101001: color_data = 12'b001110100111;
		16'b1001000010101010: color_data = 12'b001110100111;
		16'b1001000010101011: color_data = 12'b001110100111;
		16'b1001000010111000: color_data = 12'b001110100111;
		16'b1001000010111001: color_data = 12'b001110100111;
		16'b1001000010111010: color_data = 12'b001110100111;
		16'b1001000010111011: color_data = 12'b001110100111;
		16'b1001000010111100: color_data = 12'b001110100111;
		16'b1001000010111101: color_data = 12'b001110100111;
		16'b1001000010111110: color_data = 12'b001110100111;
		16'b1001000010111111: color_data = 12'b001110100111;
		16'b1001000011000000: color_data = 12'b001110100111;
		16'b1001000011000001: color_data = 12'b001110100111;
		16'b1001000011000010: color_data = 12'b001110100111;
		16'b1001000011000011: color_data = 12'b001110100111;
		16'b1001000011000100: color_data = 12'b001110100111;
		16'b1001000011001011: color_data = 12'b001110100111;
		16'b1001000011001100: color_data = 12'b001110100111;
		16'b1001000011001101: color_data = 12'b001110100111;
		16'b1001000011001110: color_data = 12'b001110100111;
		16'b1001000011001111: color_data = 12'b001110100111;
		16'b1001000011010000: color_data = 12'b001110100111;
		16'b1001000011010001: color_data = 12'b001110100111;
		16'b1001000011010010: color_data = 12'b001110100111;
		16'b1001000011010011: color_data = 12'b001110100111;
		16'b1001000011010100: color_data = 12'b001110100111;
		16'b1001000011010101: color_data = 12'b001110100111;
		16'b1001000011010110: color_data = 12'b001110100111;
		16'b1001000011110110: color_data = 12'b001110100111;
		16'b1001000011110111: color_data = 12'b001110100111;
		16'b1001000011111000: color_data = 12'b001110100111;
		16'b1001000011111001: color_data = 12'b001110100111;
		16'b1001000011111010: color_data = 12'b001110100111;
		16'b1001000011111011: color_data = 12'b001110100111;
		16'b1001000011111100: color_data = 12'b001110100111;
		16'b1001000011111101: color_data = 12'b001110100111;
		16'b1001000011111110: color_data = 12'b001110100111;
		16'b1001000011111111: color_data = 12'b001110100111;
		16'b1001000100000000: color_data = 12'b001110100111;
		16'b1001000100000001: color_data = 12'b001110100111;
		16'b1001000100011010: color_data = 12'b001110100111;
		16'b1001000100011011: color_data = 12'b001110100111;
		16'b1001000100011100: color_data = 12'b001110100111;
		16'b1001000100011101: color_data = 12'b001110100111;
		16'b1001000100011110: color_data = 12'b001110100111;
		16'b1001000100011111: color_data = 12'b001110100111;
		16'b1001000100100000: color_data = 12'b001110100111;
		16'b1001000100100001: color_data = 12'b001110100111;
		16'b1001000100100010: color_data = 12'b001110100111;
		16'b1001000100100011: color_data = 12'b001110100111;
		16'b1001000100100100: color_data = 12'b001110100111;
		16'b1001000100100101: color_data = 12'b001110100111;
		16'b1001000100100110: color_data = 12'b001110100111;
		16'b1001000100101101: color_data = 12'b001110100111;
		16'b1001000100101110: color_data = 12'b001110100111;
		16'b1001000100101111: color_data = 12'b001110100111;
		16'b1001000100110000: color_data = 12'b001110100111;
		16'b1001000100110001: color_data = 12'b001110100111;
		16'b1001000100110010: color_data = 12'b001110100111;
		16'b1001000100110011: color_data = 12'b001110100111;
		16'b1001000100110100: color_data = 12'b001110100111;
		16'b1001000100110101: color_data = 12'b001110100111;
		16'b1001000100110110: color_data = 12'b001110100111;
		16'b1001000100110111: color_data = 12'b001110100111;
		16'b1001000100111000: color_data = 12'b001110100111;
		16'b1001000101000101: color_data = 12'b001110100111;
		16'b1001000101000110: color_data = 12'b001110100111;
		16'b1001000101000111: color_data = 12'b001110100111;
		16'b1001000101001000: color_data = 12'b001110100111;
		16'b1001000101001001: color_data = 12'b001110100111;
		16'b1001000101001010: color_data = 12'b001110100111;
		16'b1001000101001011: color_data = 12'b001110100111;
		16'b1001000101001100: color_data = 12'b001110100111;
		16'b1001000101001101: color_data = 12'b001110100111;
		16'b1001000101001110: color_data = 12'b001110100111;
		16'b1001000101001111: color_data = 12'b001110100111;
		16'b1001000101010000: color_data = 12'b001110100111;
		16'b1001000101010001: color_data = 12'b001110100111;
		16'b1001000101011000: color_data = 12'b001110100111;
		16'b1001000101011001: color_data = 12'b001110100111;
		16'b1001000101011010: color_data = 12'b001110100111;
		16'b1001000101011011: color_data = 12'b001110100111;
		16'b1001000101011100: color_data = 12'b001110100111;
		16'b1001000101011101: color_data = 12'b001110100111;
		16'b1001000101011110: color_data = 12'b001110100111;
		16'b1001000101011111: color_data = 12'b001110100111;
		16'b1001000101100000: color_data = 12'b001110100111;
		16'b1001000101100001: color_data = 12'b001110100111;
		16'b1001000101100010: color_data = 12'b001110100111;
		16'b1001000101100011: color_data = 12'b001110100111;
		16'b1001000101110000: color_data = 12'b001110100111;
		16'b1001000101110001: color_data = 12'b001110100111;
		16'b1001000101110010: color_data = 12'b001110100111;
		16'b1001000101110011: color_data = 12'b001110100111;
		16'b1001000101110100: color_data = 12'b001110100111;
		16'b1001000101110101: color_data = 12'b001110100111;
		16'b1001000101110110: color_data = 12'b001110100111;
		16'b1001000101110111: color_data = 12'b001110100111;
		16'b1001000101111000: color_data = 12'b001110100111;
		16'b1001000101111001: color_data = 12'b001110100111;
		16'b1001000101111010: color_data = 12'b001110100111;
		16'b1001000101111011: color_data = 12'b001110100111;
		16'b1001001000000000: color_data = 12'b001110100111;
		16'b1001001000000001: color_data = 12'b001110100111;
		16'b1001001000000010: color_data = 12'b001110100111;
		16'b1001001000000011: color_data = 12'b001110100111;
		16'b1001001000000100: color_data = 12'b001110100111;
		16'b1001001000000101: color_data = 12'b001110100111;
		16'b1001001000000110: color_data = 12'b001110100111;
		16'b1001001000000111: color_data = 12'b001110100111;
		16'b1001001000001000: color_data = 12'b001110100111;
		16'b1001001000001001: color_data = 12'b001110100111;
		16'b1001001000001010: color_data = 12'b001110100111;
		16'b1001001000001011: color_data = 12'b001110100111;
		16'b1001001000001100: color_data = 12'b001110100111;
		16'b1001001000101011: color_data = 12'b001110100111;
		16'b1001001000101100: color_data = 12'b001110100111;
		16'b1001001000101101: color_data = 12'b001110100111;
		16'b1001001000101110: color_data = 12'b001110100111;
		16'b1001001000101111: color_data = 12'b001110100111;
		16'b1001001000110000: color_data = 12'b001110100111;
		16'b1001001000110001: color_data = 12'b001110100111;
		16'b1001001000110010: color_data = 12'b001110100111;
		16'b1001001000110011: color_data = 12'b001110100111;
		16'b1001001000110100: color_data = 12'b001110100111;
		16'b1001001000110101: color_data = 12'b001110100111;
		16'b1001001000110110: color_data = 12'b001110100111;
		16'b1001001000110111: color_data = 12'b001110100111;
		16'b1001001001000100: color_data = 12'b001110100111;
		16'b1001001001000101: color_data = 12'b001110100111;
		16'b1001001001000110: color_data = 12'b001110100111;
		16'b1001001001000111: color_data = 12'b001110100111;
		16'b1001001001001000: color_data = 12'b001110100111;
		16'b1001001001001001: color_data = 12'b001110100111;
		16'b1001001001001010: color_data = 12'b001110100111;
		16'b1001001001001011: color_data = 12'b001110100111;
		16'b1001001001001100: color_data = 12'b001110100111;
		16'b1001001001001101: color_data = 12'b001110100111;
		16'b1001001001001110: color_data = 12'b001110100111;
		16'b1001001001001111: color_data = 12'b001110100111;
		16'b1001001001011100: color_data = 12'b001110100111;
		16'b1001001001011101: color_data = 12'b001110100111;
		16'b1001001001011110: color_data = 12'b001110100111;
		16'b1001001001011111: color_data = 12'b001110100111;
		16'b1001001001100000: color_data = 12'b001110100111;
		16'b1001001001100001: color_data = 12'b001110100111;
		16'b1001001001100010: color_data = 12'b001110100111;
		16'b1001001001100011: color_data = 12'b001110100111;
		16'b1001001001100100: color_data = 12'b001110100111;
		16'b1001001001100101: color_data = 12'b001110100111;
		16'b1001001001100110: color_data = 12'b001110100111;
		16'b1001001001100111: color_data = 12'b001110100111;
		16'b1001001001101000: color_data = 12'b001110100111;
		16'b1001001001110101: color_data = 12'b001110100111;
		16'b1001001001110110: color_data = 12'b001110100111;
		16'b1001001001110111: color_data = 12'b001110100111;
		16'b1001001001111000: color_data = 12'b001110100111;
		16'b1001001001111001: color_data = 12'b001110100111;
		16'b1001001001111010: color_data = 12'b001110100111;
		16'b1001001001111011: color_data = 12'b001110100111;
		16'b1001001001111100: color_data = 12'b001110100111;
		16'b1001001001111101: color_data = 12'b001110100111;
		16'b1001001001111110: color_data = 12'b001110100111;
		16'b1001001001111111: color_data = 12'b001110100111;
		16'b1001001010000000: color_data = 12'b001110100111;
		16'b1001001010001101: color_data = 12'b001110100111;
		16'b1001001010001110: color_data = 12'b001110100111;
		16'b1001001010001111: color_data = 12'b001110100111;
		16'b1001001010010000: color_data = 12'b001110100111;
		16'b1001001010010001: color_data = 12'b001110100111;
		16'b1001001010010010: color_data = 12'b001110100111;
		16'b1001001010010011: color_data = 12'b001110100111;
		16'b1001001010010100: color_data = 12'b001110100111;
		16'b1001001010010101: color_data = 12'b001110100111;
		16'b1001001010010110: color_data = 12'b001110100111;
		16'b1001001010010111: color_data = 12'b001110100111;
		16'b1001001010011000: color_data = 12'b001110100111;
		16'b1001001010011001: color_data = 12'b001110100111;
		16'b1001001010100000: color_data = 12'b001110100111;
		16'b1001001010100001: color_data = 12'b001110100111;
		16'b1001001010100010: color_data = 12'b001110100111;
		16'b1001001010100011: color_data = 12'b001110100111;
		16'b1001001010100100: color_data = 12'b001110100111;
		16'b1001001010100101: color_data = 12'b001110100111;
		16'b1001001010100110: color_data = 12'b001110100111;
		16'b1001001010100111: color_data = 12'b001110100111;
		16'b1001001010101000: color_data = 12'b001110100111;
		16'b1001001010101001: color_data = 12'b001110100111;
		16'b1001001010101010: color_data = 12'b001110100111;
		16'b1001001010101011: color_data = 12'b001110100111;
		16'b1001001010111000: color_data = 12'b001110100111;
		16'b1001001010111001: color_data = 12'b001110100111;
		16'b1001001010111010: color_data = 12'b001110100111;
		16'b1001001010111011: color_data = 12'b001110100111;
		16'b1001001010111100: color_data = 12'b001110100111;
		16'b1001001010111101: color_data = 12'b001110100111;
		16'b1001001010111110: color_data = 12'b001110100111;
		16'b1001001010111111: color_data = 12'b001110100111;
		16'b1001001011000000: color_data = 12'b001110100111;
		16'b1001001011000001: color_data = 12'b001110100111;
		16'b1001001011000010: color_data = 12'b001110100111;
		16'b1001001011000011: color_data = 12'b001110100111;
		16'b1001001011000100: color_data = 12'b001110100111;
		16'b1001001011001011: color_data = 12'b001110100111;
		16'b1001001011001100: color_data = 12'b001110100111;
		16'b1001001011001101: color_data = 12'b001110100111;
		16'b1001001011001110: color_data = 12'b001110100111;
		16'b1001001011001111: color_data = 12'b001110100111;
		16'b1001001011010000: color_data = 12'b001110100111;
		16'b1001001011010001: color_data = 12'b001110100111;
		16'b1001001011010010: color_data = 12'b001110100111;
		16'b1001001011010011: color_data = 12'b001110100111;
		16'b1001001011010100: color_data = 12'b001110100111;
		16'b1001001011010101: color_data = 12'b001110100111;
		16'b1001001011010110: color_data = 12'b001110100111;
		16'b1001001011110110: color_data = 12'b001110100111;
		16'b1001001011110111: color_data = 12'b001110100111;
		16'b1001001011111000: color_data = 12'b001110100111;
		16'b1001001011111001: color_data = 12'b001110100111;
		16'b1001001011111010: color_data = 12'b001110100111;
		16'b1001001011111011: color_data = 12'b001110100111;
		16'b1001001011111100: color_data = 12'b001110100111;
		16'b1001001011111101: color_data = 12'b001110100111;
		16'b1001001011111110: color_data = 12'b001110100111;
		16'b1001001011111111: color_data = 12'b001110100111;
		16'b1001001100000000: color_data = 12'b001110100111;
		16'b1001001100000001: color_data = 12'b001110100111;
		16'b1001001100011010: color_data = 12'b001110100111;
		16'b1001001100011011: color_data = 12'b001110100111;
		16'b1001001100011100: color_data = 12'b001110100111;
		16'b1001001100011101: color_data = 12'b001110100111;
		16'b1001001100011110: color_data = 12'b001110100111;
		16'b1001001100011111: color_data = 12'b001110100111;
		16'b1001001100100000: color_data = 12'b001110100111;
		16'b1001001100100001: color_data = 12'b001110100111;
		16'b1001001100100010: color_data = 12'b001110100111;
		16'b1001001100100011: color_data = 12'b001110100111;
		16'b1001001100100100: color_data = 12'b001110100111;
		16'b1001001100100101: color_data = 12'b001110100111;
		16'b1001001100100110: color_data = 12'b001110100111;
		16'b1001001100101101: color_data = 12'b001110100111;
		16'b1001001100101110: color_data = 12'b001110100111;
		16'b1001001100101111: color_data = 12'b001110100111;
		16'b1001001100110000: color_data = 12'b001110100111;
		16'b1001001100110001: color_data = 12'b001110100111;
		16'b1001001100110010: color_data = 12'b001110100111;
		16'b1001001100110011: color_data = 12'b001110100111;
		16'b1001001100110100: color_data = 12'b001110100111;
		16'b1001001100110101: color_data = 12'b001110100111;
		16'b1001001100110110: color_data = 12'b001110100111;
		16'b1001001100110111: color_data = 12'b001110100111;
		16'b1001001100111000: color_data = 12'b001110100111;
		16'b1001001101000101: color_data = 12'b001110100111;
		16'b1001001101000110: color_data = 12'b001110100111;
		16'b1001001101000111: color_data = 12'b001110100111;
		16'b1001001101001000: color_data = 12'b001110100111;
		16'b1001001101001001: color_data = 12'b001110100111;
		16'b1001001101001010: color_data = 12'b001110100111;
		16'b1001001101001011: color_data = 12'b001110100111;
		16'b1001001101001100: color_data = 12'b001110100111;
		16'b1001001101001101: color_data = 12'b001110100111;
		16'b1001001101001110: color_data = 12'b001110100111;
		16'b1001001101001111: color_data = 12'b001110100111;
		16'b1001001101010000: color_data = 12'b001110100111;
		16'b1001001101010001: color_data = 12'b001110100111;
		16'b1001001101011000: color_data = 12'b001110100111;
		16'b1001001101011001: color_data = 12'b001110100111;
		16'b1001001101011010: color_data = 12'b001110100111;
		16'b1001001101011011: color_data = 12'b001110100111;
		16'b1001001101011100: color_data = 12'b001110100111;
		16'b1001001101011101: color_data = 12'b001110100111;
		16'b1001001101011110: color_data = 12'b001110100111;
		16'b1001001101011111: color_data = 12'b001110100111;
		16'b1001001101100000: color_data = 12'b001110100111;
		16'b1001001101100001: color_data = 12'b001110100111;
		16'b1001001101100010: color_data = 12'b001110100111;
		16'b1001001101100011: color_data = 12'b001110100111;
		16'b1001001101110000: color_data = 12'b001110100111;
		16'b1001001101110001: color_data = 12'b001110100111;
		16'b1001001101110010: color_data = 12'b001110100111;
		16'b1001001101110011: color_data = 12'b001110100111;
		16'b1001001101110100: color_data = 12'b001110100111;
		16'b1001001101110101: color_data = 12'b001110100111;
		16'b1001001101110110: color_data = 12'b001110100111;
		16'b1001001101110111: color_data = 12'b001110100111;
		16'b1001001101111000: color_data = 12'b001110100111;
		16'b1001001101111001: color_data = 12'b001110100111;
		16'b1001001101111010: color_data = 12'b001110100111;
		16'b1001001101111011: color_data = 12'b001110100111;
		16'b1001010000000000: color_data = 12'b001110100111;
		16'b1001010000000001: color_data = 12'b001110100111;
		16'b1001010000000010: color_data = 12'b001110100111;
		16'b1001010000000011: color_data = 12'b001110100111;
		16'b1001010000000100: color_data = 12'b001110100111;
		16'b1001010000000101: color_data = 12'b001110100111;
		16'b1001010000000110: color_data = 12'b001110100111;
		16'b1001010000000111: color_data = 12'b001110100111;
		16'b1001010000001000: color_data = 12'b001110100111;
		16'b1001010000001001: color_data = 12'b001110100111;
		16'b1001010000001010: color_data = 12'b001110100111;
		16'b1001010000001011: color_data = 12'b001110100111;
		16'b1001010000001100: color_data = 12'b001110100111;
		16'b1001010000101011: color_data = 12'b001110100111;
		16'b1001010000101100: color_data = 12'b001110100111;
		16'b1001010000101101: color_data = 12'b001110100111;
		16'b1001010000101110: color_data = 12'b001110100111;
		16'b1001010000101111: color_data = 12'b001110100111;
		16'b1001010000110000: color_data = 12'b001110100111;
		16'b1001010000110001: color_data = 12'b001110100111;
		16'b1001010000110010: color_data = 12'b001110100111;
		16'b1001010000110011: color_data = 12'b001110100111;
		16'b1001010000110100: color_data = 12'b001110100111;
		16'b1001010000110101: color_data = 12'b001110100111;
		16'b1001010000110110: color_data = 12'b001110100111;
		16'b1001010000110111: color_data = 12'b001110100111;
		16'b1001010001000100: color_data = 12'b001110100111;
		16'b1001010001000101: color_data = 12'b001110100111;
		16'b1001010001000110: color_data = 12'b001110100111;
		16'b1001010001000111: color_data = 12'b001110100111;
		16'b1001010001001000: color_data = 12'b001110100111;
		16'b1001010001001001: color_data = 12'b001110100111;
		16'b1001010001001010: color_data = 12'b001110100111;
		16'b1001010001001011: color_data = 12'b001110100111;
		16'b1001010001001100: color_data = 12'b001110100111;
		16'b1001010001001101: color_data = 12'b001110100111;
		16'b1001010001001110: color_data = 12'b001110100111;
		16'b1001010001001111: color_data = 12'b001110100111;
		16'b1001010001011100: color_data = 12'b001110100111;
		16'b1001010001011101: color_data = 12'b001110100111;
		16'b1001010001011110: color_data = 12'b001110100111;
		16'b1001010001011111: color_data = 12'b001110100111;
		16'b1001010001100000: color_data = 12'b001110100111;
		16'b1001010001100001: color_data = 12'b001110100111;
		16'b1001010001100010: color_data = 12'b001110100111;
		16'b1001010001100011: color_data = 12'b001110100111;
		16'b1001010001100100: color_data = 12'b001110100111;
		16'b1001010001100101: color_data = 12'b001110100111;
		16'b1001010001100110: color_data = 12'b001110100111;
		16'b1001010001100111: color_data = 12'b001110100111;
		16'b1001010001101000: color_data = 12'b001110100111;
		16'b1001010001110101: color_data = 12'b001110100111;
		16'b1001010001110110: color_data = 12'b001110100111;
		16'b1001010001110111: color_data = 12'b001110100111;
		16'b1001010001111000: color_data = 12'b001110100111;
		16'b1001010001111001: color_data = 12'b001110100111;
		16'b1001010001111010: color_data = 12'b001110100111;
		16'b1001010001111011: color_data = 12'b001110100111;
		16'b1001010001111100: color_data = 12'b001110100111;
		16'b1001010001111101: color_data = 12'b001110100111;
		16'b1001010001111110: color_data = 12'b001110100111;
		16'b1001010001111111: color_data = 12'b001110100111;
		16'b1001010010000000: color_data = 12'b001110100111;
		16'b1001010010001101: color_data = 12'b001110100111;
		16'b1001010010001110: color_data = 12'b001110100111;
		16'b1001010010001111: color_data = 12'b001110100111;
		16'b1001010010010000: color_data = 12'b001110100111;
		16'b1001010010010001: color_data = 12'b001110100111;
		16'b1001010010010010: color_data = 12'b001110100111;
		16'b1001010010010011: color_data = 12'b001110100111;
		16'b1001010010010100: color_data = 12'b001110100111;
		16'b1001010010010101: color_data = 12'b001110100111;
		16'b1001010010010110: color_data = 12'b001110100111;
		16'b1001010010010111: color_data = 12'b001110100111;
		16'b1001010010011000: color_data = 12'b001110100111;
		16'b1001010010011001: color_data = 12'b001110100111;
		16'b1001010010100000: color_data = 12'b001110100111;
		16'b1001010010100001: color_data = 12'b001110100111;
		16'b1001010010100010: color_data = 12'b001110100111;
		16'b1001010010100011: color_data = 12'b001110100111;
		16'b1001010010100100: color_data = 12'b001110100111;
		16'b1001010010100101: color_data = 12'b001110100111;
		16'b1001010010100110: color_data = 12'b001110100111;
		16'b1001010010100111: color_data = 12'b001110100111;
		16'b1001010010101000: color_data = 12'b001110100111;
		16'b1001010010101001: color_data = 12'b001110100111;
		16'b1001010010101010: color_data = 12'b001110100111;
		16'b1001010010101011: color_data = 12'b001110100111;
		16'b1001010010111000: color_data = 12'b001110100111;
		16'b1001010010111001: color_data = 12'b001110100111;
		16'b1001010010111010: color_data = 12'b001110100111;
		16'b1001010010111011: color_data = 12'b001110100111;
		16'b1001010010111100: color_data = 12'b001110100111;
		16'b1001010010111101: color_data = 12'b001110100111;
		16'b1001010010111110: color_data = 12'b001110100111;
		16'b1001010010111111: color_data = 12'b001110100111;
		16'b1001010011000000: color_data = 12'b001110100111;
		16'b1001010011000001: color_data = 12'b001110100111;
		16'b1001010011000010: color_data = 12'b001110100111;
		16'b1001010011000011: color_data = 12'b001110100111;
		16'b1001010011000100: color_data = 12'b001110100111;
		16'b1001010011001011: color_data = 12'b001110100111;
		16'b1001010011001100: color_data = 12'b001110100111;
		16'b1001010011001101: color_data = 12'b001110100111;
		16'b1001010011001110: color_data = 12'b001110100111;
		16'b1001010011001111: color_data = 12'b001110100111;
		16'b1001010011010000: color_data = 12'b001110100111;
		16'b1001010011010001: color_data = 12'b001110100111;
		16'b1001010011010010: color_data = 12'b001110100111;
		16'b1001010011010011: color_data = 12'b001110100111;
		16'b1001010011010100: color_data = 12'b001110100111;
		16'b1001010011010101: color_data = 12'b001110100111;
		16'b1001010011010110: color_data = 12'b001110100111;
		16'b1001010011110110: color_data = 12'b001110100111;
		16'b1001010011110111: color_data = 12'b001110100111;
		16'b1001010011111000: color_data = 12'b001110100111;
		16'b1001010011111001: color_data = 12'b001110100111;
		16'b1001010011111010: color_data = 12'b001110100111;
		16'b1001010011111011: color_data = 12'b001110100111;
		16'b1001010011111100: color_data = 12'b001110100111;
		16'b1001010011111101: color_data = 12'b001110100111;
		16'b1001010011111110: color_data = 12'b001110100111;
		16'b1001010011111111: color_data = 12'b001110100111;
		16'b1001010100000000: color_data = 12'b001110100111;
		16'b1001010100000001: color_data = 12'b001110100111;
		16'b1001010100011010: color_data = 12'b001110100111;
		16'b1001010100011011: color_data = 12'b001110100111;
		16'b1001010100011100: color_data = 12'b001110100111;
		16'b1001010100011101: color_data = 12'b001110100111;
		16'b1001010100011110: color_data = 12'b001110100111;
		16'b1001010100011111: color_data = 12'b001110100111;
		16'b1001010100100000: color_data = 12'b001110100111;
		16'b1001010100100001: color_data = 12'b001110100111;
		16'b1001010100100010: color_data = 12'b001110100111;
		16'b1001010100100011: color_data = 12'b001110100111;
		16'b1001010100100100: color_data = 12'b001110100111;
		16'b1001010100100101: color_data = 12'b001110100111;
		16'b1001010100100110: color_data = 12'b001110100111;
		16'b1001010100101101: color_data = 12'b001110100111;
		16'b1001010100101110: color_data = 12'b001110100111;
		16'b1001010100101111: color_data = 12'b001110100111;
		16'b1001010100110000: color_data = 12'b001110100111;
		16'b1001010100110001: color_data = 12'b001110100111;
		16'b1001010100110010: color_data = 12'b001110100111;
		16'b1001010100110011: color_data = 12'b001110100111;
		16'b1001010100110100: color_data = 12'b001110100111;
		16'b1001010100110101: color_data = 12'b001110100111;
		16'b1001010100110110: color_data = 12'b001110100111;
		16'b1001010100110111: color_data = 12'b001110100111;
		16'b1001010100111000: color_data = 12'b001110100111;
		16'b1001010101000101: color_data = 12'b001110100111;
		16'b1001010101000110: color_data = 12'b001110100111;
		16'b1001010101000111: color_data = 12'b001110100111;
		16'b1001010101001000: color_data = 12'b001110100111;
		16'b1001010101001001: color_data = 12'b001110100111;
		16'b1001010101001010: color_data = 12'b001110100111;
		16'b1001010101001011: color_data = 12'b001110100111;
		16'b1001010101001100: color_data = 12'b001110100111;
		16'b1001010101001101: color_data = 12'b001110100111;
		16'b1001010101001110: color_data = 12'b001110100111;
		16'b1001010101001111: color_data = 12'b001110100111;
		16'b1001010101010000: color_data = 12'b001110100111;
		16'b1001010101010001: color_data = 12'b001110100111;
		16'b1001010101011000: color_data = 12'b001110100111;
		16'b1001010101011001: color_data = 12'b001110100111;
		16'b1001010101011010: color_data = 12'b001110100111;
		16'b1001010101011011: color_data = 12'b001110100111;
		16'b1001010101011100: color_data = 12'b001110100111;
		16'b1001010101011101: color_data = 12'b001110100111;
		16'b1001010101011110: color_data = 12'b001110100111;
		16'b1001010101011111: color_data = 12'b001110100111;
		16'b1001010101100000: color_data = 12'b001110100111;
		16'b1001010101100001: color_data = 12'b001110100111;
		16'b1001010101100010: color_data = 12'b001110100111;
		16'b1001010101100011: color_data = 12'b001110100111;
		16'b1001010101110000: color_data = 12'b001110100111;
		16'b1001010101110001: color_data = 12'b001110100111;
		16'b1001010101110010: color_data = 12'b001110100111;
		16'b1001010101110011: color_data = 12'b001110100111;
		16'b1001010101110100: color_data = 12'b001110100111;
		16'b1001010101110101: color_data = 12'b001110100111;
		16'b1001010101110110: color_data = 12'b001110100111;
		16'b1001010101110111: color_data = 12'b001110100111;
		16'b1001010101111000: color_data = 12'b001110100111;
		16'b1001010101111001: color_data = 12'b001110100111;
		16'b1001010101111010: color_data = 12'b001110100111;
		16'b1001010101111011: color_data = 12'b001110100111;
		16'b1001011000000000: color_data = 12'b001110100111;
		16'b1001011000000001: color_data = 12'b001110100111;
		16'b1001011000000010: color_data = 12'b001110100111;
		16'b1001011000000011: color_data = 12'b001110100111;
		16'b1001011000000100: color_data = 12'b001110100111;
		16'b1001011000000101: color_data = 12'b001110100111;
		16'b1001011000000110: color_data = 12'b001110100111;
		16'b1001011000000111: color_data = 12'b001110100111;
		16'b1001011000001000: color_data = 12'b001110100111;
		16'b1001011000001001: color_data = 12'b001110100111;
		16'b1001011000001010: color_data = 12'b001110100111;
		16'b1001011000001011: color_data = 12'b001110100111;
		16'b1001011000001100: color_data = 12'b001110100111;
		16'b1001011000101011: color_data = 12'b001110100111;
		16'b1001011000101100: color_data = 12'b001110100111;
		16'b1001011000101101: color_data = 12'b001110100111;
		16'b1001011000101110: color_data = 12'b001110100111;
		16'b1001011000101111: color_data = 12'b001110100111;
		16'b1001011000110000: color_data = 12'b001110100111;
		16'b1001011000110001: color_data = 12'b001110100111;
		16'b1001011000110010: color_data = 12'b001110100111;
		16'b1001011000110011: color_data = 12'b001110100111;
		16'b1001011000110100: color_data = 12'b001110100111;
		16'b1001011000110101: color_data = 12'b001110100111;
		16'b1001011000110110: color_data = 12'b001110100111;
		16'b1001011000110111: color_data = 12'b001110100111;
		16'b1001011001000100: color_data = 12'b001110100111;
		16'b1001011001000101: color_data = 12'b001110100111;
		16'b1001011001000110: color_data = 12'b001110100111;
		16'b1001011001000111: color_data = 12'b001110100111;
		16'b1001011001001000: color_data = 12'b001110100111;
		16'b1001011001001001: color_data = 12'b001110100111;
		16'b1001011001001010: color_data = 12'b001110100111;
		16'b1001011001001011: color_data = 12'b001110100111;
		16'b1001011001001100: color_data = 12'b001110100111;
		16'b1001011001001101: color_data = 12'b001110100111;
		16'b1001011001001110: color_data = 12'b001110100111;
		16'b1001011001001111: color_data = 12'b001110100111;
		16'b1001011001011100: color_data = 12'b001110100111;
		16'b1001011001011101: color_data = 12'b001110100111;
		16'b1001011001011110: color_data = 12'b001110100111;
		16'b1001011001011111: color_data = 12'b001110100111;
		16'b1001011001100000: color_data = 12'b001110100111;
		16'b1001011001100001: color_data = 12'b001110100111;
		16'b1001011001100010: color_data = 12'b001110100111;
		16'b1001011001100011: color_data = 12'b001110100111;
		16'b1001011001100100: color_data = 12'b001110100111;
		16'b1001011001100101: color_data = 12'b001110100111;
		16'b1001011001100110: color_data = 12'b001110100111;
		16'b1001011001100111: color_data = 12'b001110100111;
		16'b1001011001101000: color_data = 12'b001110100111;
		16'b1001011001110101: color_data = 12'b001110100111;
		16'b1001011001110110: color_data = 12'b001110100111;
		16'b1001011001110111: color_data = 12'b001110100111;
		16'b1001011001111000: color_data = 12'b001110100111;
		16'b1001011001111001: color_data = 12'b001110100111;
		16'b1001011001111010: color_data = 12'b001110100111;
		16'b1001011001111011: color_data = 12'b001110100111;
		16'b1001011001111100: color_data = 12'b001110100111;
		16'b1001011001111101: color_data = 12'b001110100111;
		16'b1001011001111110: color_data = 12'b001110100111;
		16'b1001011001111111: color_data = 12'b001110100111;
		16'b1001011010000000: color_data = 12'b001110100111;
		16'b1001011010001101: color_data = 12'b001110100111;
		16'b1001011010001110: color_data = 12'b001110100111;
		16'b1001011010001111: color_data = 12'b001110100111;
		16'b1001011010010000: color_data = 12'b001110100111;
		16'b1001011010010001: color_data = 12'b001110100111;
		16'b1001011010010010: color_data = 12'b001110100111;
		16'b1001011010010011: color_data = 12'b001110100111;
		16'b1001011010010100: color_data = 12'b001110100111;
		16'b1001011010010101: color_data = 12'b001110100111;
		16'b1001011010010110: color_data = 12'b001110100111;
		16'b1001011010010111: color_data = 12'b001110100111;
		16'b1001011010011000: color_data = 12'b001110100111;
		16'b1001011010011001: color_data = 12'b001110100111;
		16'b1001011010100000: color_data = 12'b001110100111;
		16'b1001011010100001: color_data = 12'b001110100111;
		16'b1001011010100010: color_data = 12'b001110100111;
		16'b1001011010100011: color_data = 12'b001110100111;
		16'b1001011010100100: color_data = 12'b001110100111;
		16'b1001011010100101: color_data = 12'b001110100111;
		16'b1001011010100110: color_data = 12'b001110100111;
		16'b1001011010100111: color_data = 12'b001110100111;
		16'b1001011010101000: color_data = 12'b001110100111;
		16'b1001011010101001: color_data = 12'b001110100111;
		16'b1001011010101010: color_data = 12'b001110100111;
		16'b1001011010101011: color_data = 12'b001110100111;
		16'b1001011010111000: color_data = 12'b001110100111;
		16'b1001011010111001: color_data = 12'b001110100111;
		16'b1001011010111010: color_data = 12'b001110100111;
		16'b1001011010111011: color_data = 12'b001110100111;
		16'b1001011010111100: color_data = 12'b001110100111;
		16'b1001011010111101: color_data = 12'b001110100111;
		16'b1001011010111110: color_data = 12'b001110100111;
		16'b1001011010111111: color_data = 12'b001110100111;
		16'b1001011011000000: color_data = 12'b001110100111;
		16'b1001011011000001: color_data = 12'b001110100111;
		16'b1001011011000010: color_data = 12'b001110100111;
		16'b1001011011000011: color_data = 12'b001110100111;
		16'b1001011011000100: color_data = 12'b001110100111;
		16'b1001011011001011: color_data = 12'b001110100111;
		16'b1001011011001100: color_data = 12'b001110100111;
		16'b1001011011001101: color_data = 12'b001110100111;
		16'b1001011011001110: color_data = 12'b001110100111;
		16'b1001011011001111: color_data = 12'b001110100111;
		16'b1001011011010000: color_data = 12'b001110100111;
		16'b1001011011010001: color_data = 12'b001110100111;
		16'b1001011011010010: color_data = 12'b001110100111;
		16'b1001011011010011: color_data = 12'b001110100111;
		16'b1001011011010100: color_data = 12'b001110100111;
		16'b1001011011010101: color_data = 12'b001110100111;
		16'b1001011011010110: color_data = 12'b001110100111;
		16'b1001011011110110: color_data = 12'b001110100111;
		16'b1001011011110111: color_data = 12'b001110100111;
		16'b1001011011111000: color_data = 12'b001110100111;
		16'b1001011011111001: color_data = 12'b001110100111;
		16'b1001011011111010: color_data = 12'b001110100111;
		16'b1001011011111011: color_data = 12'b001110100111;
		16'b1001011011111100: color_data = 12'b001110100111;
		16'b1001011011111101: color_data = 12'b001110100111;
		16'b1001011011111110: color_data = 12'b001110100111;
		16'b1001011011111111: color_data = 12'b001110100111;
		16'b1001011100000000: color_data = 12'b001110100111;
		16'b1001011100000001: color_data = 12'b001110100111;
		16'b1001011100011010: color_data = 12'b001110100111;
		16'b1001011100011011: color_data = 12'b001110100111;
		16'b1001011100011100: color_data = 12'b001110100111;
		16'b1001011100011101: color_data = 12'b001110100111;
		16'b1001011100011110: color_data = 12'b001110100111;
		16'b1001011100011111: color_data = 12'b001110100111;
		16'b1001011100100000: color_data = 12'b001110100111;
		16'b1001011100100001: color_data = 12'b001110100111;
		16'b1001011100100010: color_data = 12'b001110100111;
		16'b1001011100100011: color_data = 12'b001110100111;
		16'b1001011100100100: color_data = 12'b001110100111;
		16'b1001011100100101: color_data = 12'b001110100111;
		16'b1001011100100110: color_data = 12'b001110100111;
		16'b1001011100101101: color_data = 12'b001110100111;
		16'b1001011100101110: color_data = 12'b001110100111;
		16'b1001011100101111: color_data = 12'b001110100111;
		16'b1001011100110000: color_data = 12'b001110100111;
		16'b1001011100110001: color_data = 12'b001110100111;
		16'b1001011100110010: color_data = 12'b001110100111;
		16'b1001011100110011: color_data = 12'b001110100111;
		16'b1001011100110100: color_data = 12'b001110100111;
		16'b1001011100110101: color_data = 12'b001110100111;
		16'b1001011100110110: color_data = 12'b001110100111;
		16'b1001011100110111: color_data = 12'b001110100111;
		16'b1001011100111000: color_data = 12'b001110100111;
		16'b1001011101000101: color_data = 12'b001110100111;
		16'b1001011101000110: color_data = 12'b001110100111;
		16'b1001011101000111: color_data = 12'b001110100111;
		16'b1001011101001000: color_data = 12'b001110100111;
		16'b1001011101001001: color_data = 12'b001110100111;
		16'b1001011101001010: color_data = 12'b001110100111;
		16'b1001011101001011: color_data = 12'b001110100111;
		16'b1001011101001100: color_data = 12'b001110100111;
		16'b1001011101001101: color_data = 12'b001110100111;
		16'b1001011101001110: color_data = 12'b001110100111;
		16'b1001011101001111: color_data = 12'b001110100111;
		16'b1001011101010000: color_data = 12'b001110100111;
		16'b1001011101010001: color_data = 12'b001110100111;
		16'b1001011101011000: color_data = 12'b001110100111;
		16'b1001011101011001: color_data = 12'b001110100111;
		16'b1001011101011010: color_data = 12'b001110100111;
		16'b1001011101011011: color_data = 12'b001110100111;
		16'b1001011101011100: color_data = 12'b001110100111;
		16'b1001011101011101: color_data = 12'b001110100111;
		16'b1001011101011110: color_data = 12'b001110100111;
		16'b1001011101011111: color_data = 12'b001110100111;
		16'b1001011101100000: color_data = 12'b001110100111;
		16'b1001011101100001: color_data = 12'b001110100111;
		16'b1001011101100010: color_data = 12'b001110100111;
		16'b1001011101100011: color_data = 12'b001110100111;
		16'b1001011101110000: color_data = 12'b001110100111;
		16'b1001011101110001: color_data = 12'b001110100111;
		16'b1001011101110010: color_data = 12'b001110100111;
		16'b1001011101110011: color_data = 12'b001110100111;
		16'b1001011101110100: color_data = 12'b001110100111;
		16'b1001011101110101: color_data = 12'b001110100111;
		16'b1001011101110110: color_data = 12'b001110100111;
		16'b1001011101110111: color_data = 12'b001110100111;
		16'b1001011101111000: color_data = 12'b001110100111;
		16'b1001011101111001: color_data = 12'b001110100111;
		16'b1001011101111010: color_data = 12'b001110100111;
		16'b1001011101111011: color_data = 12'b001110100111;
		16'b1001100000000000: color_data = 12'b001110100111;
		16'b1001100000000001: color_data = 12'b001110100111;
		16'b1001100000000010: color_data = 12'b001110100111;
		16'b1001100000000011: color_data = 12'b001110100111;
		16'b1001100000000100: color_data = 12'b001110100111;
		16'b1001100000000101: color_data = 12'b001110100111;
		16'b1001100000000110: color_data = 12'b001110100111;
		16'b1001100000000111: color_data = 12'b001110100111;
		16'b1001100000001000: color_data = 12'b001110100111;
		16'b1001100000001001: color_data = 12'b001110100111;
		16'b1001100000001010: color_data = 12'b001110100111;
		16'b1001100000001011: color_data = 12'b001110100111;
		16'b1001100000001100: color_data = 12'b001110100111;
		16'b1001100000101011: color_data = 12'b001110100111;
		16'b1001100000101100: color_data = 12'b001110100111;
		16'b1001100000101101: color_data = 12'b001110100111;
		16'b1001100000101110: color_data = 12'b001110100111;
		16'b1001100000101111: color_data = 12'b001110100111;
		16'b1001100000110000: color_data = 12'b001110100111;
		16'b1001100000110001: color_data = 12'b001110100111;
		16'b1001100000110010: color_data = 12'b001110100111;
		16'b1001100000110011: color_data = 12'b001110100111;
		16'b1001100000110100: color_data = 12'b001110100111;
		16'b1001100000110101: color_data = 12'b001110100111;
		16'b1001100000110110: color_data = 12'b001110100111;
		16'b1001100000110111: color_data = 12'b001110100111;
		16'b1001100001000100: color_data = 12'b001110100111;
		16'b1001100001000101: color_data = 12'b001110100111;
		16'b1001100001000110: color_data = 12'b001110100111;
		16'b1001100001000111: color_data = 12'b001110100111;
		16'b1001100001001000: color_data = 12'b001110100111;
		16'b1001100001001001: color_data = 12'b001110100111;
		16'b1001100001001010: color_data = 12'b001110100111;
		16'b1001100001001011: color_data = 12'b001110100111;
		16'b1001100001001100: color_data = 12'b001110100111;
		16'b1001100001001101: color_data = 12'b001110100111;
		16'b1001100001001110: color_data = 12'b001110100111;
		16'b1001100001001111: color_data = 12'b001110100111;
		16'b1001100001011100: color_data = 12'b001110100111;
		16'b1001100001011101: color_data = 12'b001110100111;
		16'b1001100001011110: color_data = 12'b001110100111;
		16'b1001100001011111: color_data = 12'b001110100111;
		16'b1001100001100000: color_data = 12'b001110100111;
		16'b1001100001100001: color_data = 12'b001110100111;
		16'b1001100001100010: color_data = 12'b001110100111;
		16'b1001100001100011: color_data = 12'b001110100111;
		16'b1001100001100100: color_data = 12'b001110100111;
		16'b1001100001100101: color_data = 12'b001110100111;
		16'b1001100001100110: color_data = 12'b001110100111;
		16'b1001100001100111: color_data = 12'b001110100111;
		16'b1001100001101000: color_data = 12'b001110100111;
		16'b1001100001110101: color_data = 12'b001110100111;
		16'b1001100001110110: color_data = 12'b001110100111;
		16'b1001100001110111: color_data = 12'b001110100111;
		16'b1001100001111000: color_data = 12'b001110100111;
		16'b1001100001111001: color_data = 12'b001110100111;
		16'b1001100001111010: color_data = 12'b001110100111;
		16'b1001100001111011: color_data = 12'b001110100111;
		16'b1001100001111100: color_data = 12'b001110100111;
		16'b1001100001111101: color_data = 12'b001110100111;
		16'b1001100001111110: color_data = 12'b001110100111;
		16'b1001100001111111: color_data = 12'b001110100111;
		16'b1001100010000000: color_data = 12'b001110100111;
		16'b1001100010001101: color_data = 12'b001110100111;
		16'b1001100010001110: color_data = 12'b001110100111;
		16'b1001100010001111: color_data = 12'b001110100111;
		16'b1001100010010000: color_data = 12'b001110100111;
		16'b1001100010010001: color_data = 12'b001110100111;
		16'b1001100010010010: color_data = 12'b001110100111;
		16'b1001100010010011: color_data = 12'b001110100111;
		16'b1001100010010100: color_data = 12'b001110100111;
		16'b1001100010010101: color_data = 12'b001110100111;
		16'b1001100010010110: color_data = 12'b001110100111;
		16'b1001100010010111: color_data = 12'b001110100111;
		16'b1001100010011000: color_data = 12'b001110100111;
		16'b1001100010011001: color_data = 12'b001110100111;
		16'b1001100010100000: color_data = 12'b001110100111;
		16'b1001100010100001: color_data = 12'b001110100111;
		16'b1001100010100010: color_data = 12'b001110100111;
		16'b1001100010100011: color_data = 12'b001110100111;
		16'b1001100010100100: color_data = 12'b001110100111;
		16'b1001100010100101: color_data = 12'b001110100111;
		16'b1001100010100110: color_data = 12'b001110100111;
		16'b1001100010100111: color_data = 12'b001110100111;
		16'b1001100010101000: color_data = 12'b001110100111;
		16'b1001100010101001: color_data = 12'b001110100111;
		16'b1001100010101010: color_data = 12'b001110100111;
		16'b1001100010101011: color_data = 12'b001110100111;
		16'b1001100010111000: color_data = 12'b001110100111;
		16'b1001100010111001: color_data = 12'b001110100111;
		16'b1001100010111010: color_data = 12'b001110100111;
		16'b1001100010111011: color_data = 12'b001110100111;
		16'b1001100010111100: color_data = 12'b001110100111;
		16'b1001100010111101: color_data = 12'b001110100111;
		16'b1001100010111110: color_data = 12'b001110100111;
		16'b1001100010111111: color_data = 12'b001110100111;
		16'b1001100011000000: color_data = 12'b001110100111;
		16'b1001100011000001: color_data = 12'b001110100111;
		16'b1001100011000010: color_data = 12'b001110100111;
		16'b1001100011000011: color_data = 12'b001110100111;
		16'b1001100011000100: color_data = 12'b001110100111;
		16'b1001100011001011: color_data = 12'b001110100111;
		16'b1001100011001100: color_data = 12'b001110100111;
		16'b1001100011001101: color_data = 12'b001110100111;
		16'b1001100011001110: color_data = 12'b001110100111;
		16'b1001100011001111: color_data = 12'b001110100111;
		16'b1001100011010000: color_data = 12'b001110100111;
		16'b1001100011010001: color_data = 12'b001110100111;
		16'b1001100011010010: color_data = 12'b001110100111;
		16'b1001100011010011: color_data = 12'b001110100111;
		16'b1001100011010100: color_data = 12'b001110100111;
		16'b1001100011010101: color_data = 12'b001110100111;
		16'b1001100011010110: color_data = 12'b001110100111;
		16'b1001100011110110: color_data = 12'b001110100111;
		16'b1001100011110111: color_data = 12'b001110100111;
		16'b1001100011111000: color_data = 12'b001110100111;
		16'b1001100011111001: color_data = 12'b001110100111;
		16'b1001100011111010: color_data = 12'b001110100111;
		16'b1001100011111011: color_data = 12'b001110100111;
		16'b1001100011111100: color_data = 12'b001110100111;
		16'b1001100011111101: color_data = 12'b001110100111;
		16'b1001100011111110: color_data = 12'b001110100111;
		16'b1001100011111111: color_data = 12'b001110100111;
		16'b1001100100000000: color_data = 12'b001110100111;
		16'b1001100100000001: color_data = 12'b001110100111;
		16'b1001100100011010: color_data = 12'b001110100111;
		16'b1001100100011011: color_data = 12'b001110100111;
		16'b1001100100011100: color_data = 12'b001110100111;
		16'b1001100100011101: color_data = 12'b001110100111;
		16'b1001100100011110: color_data = 12'b001110100111;
		16'b1001100100011111: color_data = 12'b001110100111;
		16'b1001100100100000: color_data = 12'b001110100111;
		16'b1001100100100001: color_data = 12'b001110100111;
		16'b1001100100100010: color_data = 12'b001110100111;
		16'b1001100100100011: color_data = 12'b001110100111;
		16'b1001100100100100: color_data = 12'b001110100111;
		16'b1001100100100101: color_data = 12'b001110100111;
		16'b1001100100100110: color_data = 12'b001110100111;
		16'b1001100100101101: color_data = 12'b001110100111;
		16'b1001100100101110: color_data = 12'b001110100111;
		16'b1001100100101111: color_data = 12'b001110100111;
		16'b1001100100110000: color_data = 12'b001110100111;
		16'b1001100100110001: color_data = 12'b001110100111;
		16'b1001100100110010: color_data = 12'b001110100111;
		16'b1001100100110011: color_data = 12'b001110100111;
		16'b1001100100110100: color_data = 12'b001110100111;
		16'b1001100100110101: color_data = 12'b001110100111;
		16'b1001100100110110: color_data = 12'b001110100111;
		16'b1001100100110111: color_data = 12'b001110100111;
		16'b1001100100111000: color_data = 12'b001110100111;
		16'b1001100101000101: color_data = 12'b001110100111;
		16'b1001100101000110: color_data = 12'b001110100111;
		16'b1001100101000111: color_data = 12'b001110100111;
		16'b1001100101001000: color_data = 12'b001110100111;
		16'b1001100101001001: color_data = 12'b001110100111;
		16'b1001100101001010: color_data = 12'b001110100111;
		16'b1001100101001011: color_data = 12'b001110100111;
		16'b1001100101001100: color_data = 12'b001110100111;
		16'b1001100101001101: color_data = 12'b001110100111;
		16'b1001100101001110: color_data = 12'b001110100111;
		16'b1001100101001111: color_data = 12'b001110100111;
		16'b1001100101010000: color_data = 12'b001110100111;
		16'b1001100101010001: color_data = 12'b001110100111;
		16'b1001100101011000: color_data = 12'b001110100111;
		16'b1001100101011001: color_data = 12'b001110100111;
		16'b1001100101011010: color_data = 12'b001110100111;
		16'b1001100101011011: color_data = 12'b001110100111;
		16'b1001100101011100: color_data = 12'b001110100111;
		16'b1001100101011101: color_data = 12'b001110100111;
		16'b1001100101011110: color_data = 12'b001110100111;
		16'b1001100101011111: color_data = 12'b001110100111;
		16'b1001100101100000: color_data = 12'b001110100111;
		16'b1001100101100001: color_data = 12'b001110100111;
		16'b1001100101100010: color_data = 12'b001110100111;
		16'b1001100101100011: color_data = 12'b001110100111;
		16'b1001100101110000: color_data = 12'b001110100111;
		16'b1001100101110001: color_data = 12'b001110100111;
		16'b1001100101110010: color_data = 12'b001110100111;
		16'b1001100101110011: color_data = 12'b001110100111;
		16'b1001100101110100: color_data = 12'b001110100111;
		16'b1001100101110101: color_data = 12'b001110100111;
		16'b1001100101110110: color_data = 12'b001110100111;
		16'b1001100101110111: color_data = 12'b001110100111;
		16'b1001100101111000: color_data = 12'b001110100111;
		16'b1001100101111001: color_data = 12'b001110100111;
		16'b1001100101111010: color_data = 12'b001110100111;
		16'b1001100101111011: color_data = 12'b001110100111;
		16'b1001101000000000: color_data = 12'b001110100111;
		16'b1001101000000001: color_data = 12'b001110100111;
		16'b1001101000000010: color_data = 12'b001110100111;
		16'b1001101000000011: color_data = 12'b001110100111;
		16'b1001101000000100: color_data = 12'b001110100111;
		16'b1001101000000101: color_data = 12'b001110100111;
		16'b1001101000000110: color_data = 12'b001110100111;
		16'b1001101000000111: color_data = 12'b001110100111;
		16'b1001101000001000: color_data = 12'b001110100111;
		16'b1001101000001001: color_data = 12'b001110100111;
		16'b1001101000001010: color_data = 12'b001110100111;
		16'b1001101000001011: color_data = 12'b001110100111;
		16'b1001101000001100: color_data = 12'b001110100111;
		16'b1001101000001101: color_data = 12'b001110100111;
		16'b1001101000001110: color_data = 12'b001110100111;
		16'b1001101000001111: color_data = 12'b001110100111;
		16'b1001101000010000: color_data = 12'b001110100111;
		16'b1001101000010001: color_data = 12'b001110100111;
		16'b1001101000010010: color_data = 12'b001110100111;
		16'b1001101000010011: color_data = 12'b001110100111;
		16'b1001101000010100: color_data = 12'b001110100111;
		16'b1001101000010101: color_data = 12'b001110100111;
		16'b1001101000010110: color_data = 12'b001110100111;
		16'b1001101000010111: color_data = 12'b001110100111;
		16'b1001101000011000: color_data = 12'b001110100111;
		16'b1001101000011001: color_data = 12'b001110100111;
		16'b1001101000011010: color_data = 12'b001110100111;
		16'b1001101000011011: color_data = 12'b001110100111;
		16'b1001101000011100: color_data = 12'b001110100111;
		16'b1001101000011101: color_data = 12'b001110100111;
		16'b1001101000011110: color_data = 12'b001110100111;
		16'b1001101000011111: color_data = 12'b001110100111;
		16'b1001101000100000: color_data = 12'b001110100111;
		16'b1001101000100001: color_data = 12'b001110100111;
		16'b1001101000100010: color_data = 12'b001110100111;
		16'b1001101000100011: color_data = 12'b001110100111;
		16'b1001101000100100: color_data = 12'b001110100111;
		16'b1001101000101011: color_data = 12'b001110100111;
		16'b1001101000101100: color_data = 12'b001110100111;
		16'b1001101000101101: color_data = 12'b001110100111;
		16'b1001101000101110: color_data = 12'b001110100111;
		16'b1001101000101111: color_data = 12'b001110100111;
		16'b1001101000110000: color_data = 12'b001110100111;
		16'b1001101000110001: color_data = 12'b001110100111;
		16'b1001101000110010: color_data = 12'b001110100111;
		16'b1001101000110011: color_data = 12'b001110100111;
		16'b1001101000110100: color_data = 12'b001110100111;
		16'b1001101000110101: color_data = 12'b001110100111;
		16'b1001101000110110: color_data = 12'b001110100111;
		16'b1001101000110111: color_data = 12'b001110100111;
		16'b1001101001000100: color_data = 12'b001110100111;
		16'b1001101001000101: color_data = 12'b001110100111;
		16'b1001101001000110: color_data = 12'b001110100111;
		16'b1001101001000111: color_data = 12'b001110100111;
		16'b1001101001001000: color_data = 12'b001110100111;
		16'b1001101001001001: color_data = 12'b001110100111;
		16'b1001101001001010: color_data = 12'b001110100111;
		16'b1001101001001011: color_data = 12'b001110100111;
		16'b1001101001001100: color_data = 12'b001110100111;
		16'b1001101001001101: color_data = 12'b001110100111;
		16'b1001101001001110: color_data = 12'b001110100111;
		16'b1001101001001111: color_data = 12'b001110100111;
		16'b1001101001010110: color_data = 12'b001110100111;
		16'b1001101001010111: color_data = 12'b001110100111;
		16'b1001101001011000: color_data = 12'b001110100111;
		16'b1001101001011001: color_data = 12'b001110100111;
		16'b1001101001011010: color_data = 12'b001110100111;
		16'b1001101001011011: color_data = 12'b001110100111;
		16'b1001101001011100: color_data = 12'b001110100111;
		16'b1001101001011101: color_data = 12'b001110100111;
		16'b1001101001011110: color_data = 12'b001110100111;
		16'b1001101001011111: color_data = 12'b001110100111;
		16'b1001101001100000: color_data = 12'b001110100111;
		16'b1001101001100001: color_data = 12'b001110100111;
		16'b1001101001100010: color_data = 12'b001110100111;
		16'b1001101001100011: color_data = 12'b001110100111;
		16'b1001101001100100: color_data = 12'b001110100111;
		16'b1001101001100101: color_data = 12'b001110100111;
		16'b1001101001100110: color_data = 12'b001110100111;
		16'b1001101001100111: color_data = 12'b001110100111;
		16'b1001101001101000: color_data = 12'b001110100111;
		16'b1001101001101001: color_data = 12'b001110100111;
		16'b1001101001101010: color_data = 12'b001110100111;
		16'b1001101001101011: color_data = 12'b001110100111;
		16'b1001101001101100: color_data = 12'b001110100111;
		16'b1001101001101101: color_data = 12'b001110100111;
		16'b1001101001101110: color_data = 12'b001110100111;
		16'b1001101001110101: color_data = 12'b001110100111;
		16'b1001101001110110: color_data = 12'b001110100111;
		16'b1001101001110111: color_data = 12'b001110100111;
		16'b1001101001111000: color_data = 12'b001110100111;
		16'b1001101001111001: color_data = 12'b001110100111;
		16'b1001101001111010: color_data = 12'b001110100111;
		16'b1001101001111011: color_data = 12'b001110100111;
		16'b1001101001111100: color_data = 12'b001110100111;
		16'b1001101001111101: color_data = 12'b001110100111;
		16'b1001101001111110: color_data = 12'b001110100111;
		16'b1001101001111111: color_data = 12'b001110100111;
		16'b1001101010000000: color_data = 12'b001110100111;
		16'b1001101010001101: color_data = 12'b001110100111;
		16'b1001101010001110: color_data = 12'b001110100111;
		16'b1001101010001111: color_data = 12'b001110100111;
		16'b1001101010010000: color_data = 12'b001110100111;
		16'b1001101010010001: color_data = 12'b001110100111;
		16'b1001101010010010: color_data = 12'b001110100111;
		16'b1001101010010011: color_data = 12'b001110100111;
		16'b1001101010010100: color_data = 12'b001110100111;
		16'b1001101010010101: color_data = 12'b001110100111;
		16'b1001101010010110: color_data = 12'b001110100111;
		16'b1001101010010111: color_data = 12'b001110100111;
		16'b1001101010011000: color_data = 12'b001110100111;
		16'b1001101010011001: color_data = 12'b001110100111;
		16'b1001101010100000: color_data = 12'b001110100111;
		16'b1001101010100001: color_data = 12'b001110100111;
		16'b1001101010100010: color_data = 12'b001110100111;
		16'b1001101010100011: color_data = 12'b001110100111;
		16'b1001101010100100: color_data = 12'b001110100111;
		16'b1001101010100101: color_data = 12'b001110100111;
		16'b1001101010100110: color_data = 12'b001110100111;
		16'b1001101010100111: color_data = 12'b001110100111;
		16'b1001101010101000: color_data = 12'b001110100111;
		16'b1001101010101001: color_data = 12'b001110100111;
		16'b1001101010101010: color_data = 12'b001110100111;
		16'b1001101010101011: color_data = 12'b001110100111;
		16'b1001101010101100: color_data = 12'b001110100111;
		16'b1001101010101101: color_data = 12'b001110100111;
		16'b1001101010101110: color_data = 12'b001110100111;
		16'b1001101010101111: color_data = 12'b001110100111;
		16'b1001101010110000: color_data = 12'b001110100111;
		16'b1001101010110001: color_data = 12'b001110100111;
		16'b1001101010110010: color_data = 12'b001110100111;
		16'b1001101010110011: color_data = 12'b001110100111;
		16'b1001101010110100: color_data = 12'b001110100111;
		16'b1001101010110101: color_data = 12'b001110100111;
		16'b1001101010110110: color_data = 12'b001110100111;
		16'b1001101010110111: color_data = 12'b001110100111;
		16'b1001101010111000: color_data = 12'b001110100111;
		16'b1001101010111001: color_data = 12'b001110100111;
		16'b1001101010111010: color_data = 12'b001110100111;
		16'b1001101010111011: color_data = 12'b001110100111;
		16'b1001101010111100: color_data = 12'b001110100111;
		16'b1001101010111101: color_data = 12'b001110100111;
		16'b1001101010111110: color_data = 12'b001110100111;
		16'b1001101010111111: color_data = 12'b001110100111;
		16'b1001101011000000: color_data = 12'b001110100111;
		16'b1001101011000001: color_data = 12'b001110100111;
		16'b1001101011000010: color_data = 12'b001110100111;
		16'b1001101011000011: color_data = 12'b001110100111;
		16'b1001101011000100: color_data = 12'b001110100111;
		16'b1001101011001011: color_data = 12'b001110100111;
		16'b1001101011001100: color_data = 12'b001110100111;
		16'b1001101011001101: color_data = 12'b001110100111;
		16'b1001101011001110: color_data = 12'b001110100111;
		16'b1001101011001111: color_data = 12'b001110100111;
		16'b1001101011010000: color_data = 12'b001110100111;
		16'b1001101011010001: color_data = 12'b001110100111;
		16'b1001101011010010: color_data = 12'b001110100111;
		16'b1001101011010011: color_data = 12'b001110100111;
		16'b1001101011010100: color_data = 12'b001110100111;
		16'b1001101011010101: color_data = 12'b001110100111;
		16'b1001101011010110: color_data = 12'b001110100111;
		16'b1001101011110110: color_data = 12'b001110100111;
		16'b1001101011110111: color_data = 12'b001110100111;
		16'b1001101011111000: color_data = 12'b001110100111;
		16'b1001101011111001: color_data = 12'b001110100111;
		16'b1001101011111010: color_data = 12'b001110100111;
		16'b1001101011111011: color_data = 12'b001110100111;
		16'b1001101011111100: color_data = 12'b001110100111;
		16'b1001101011111101: color_data = 12'b001110100111;
		16'b1001101011111110: color_data = 12'b001110100111;
		16'b1001101011111111: color_data = 12'b001110100111;
		16'b1001101100000000: color_data = 12'b001110100111;
		16'b1001101100000001: color_data = 12'b001110100111;
		16'b1001101100000010: color_data = 12'b001110100111;
		16'b1001101100000011: color_data = 12'b001110100111;
		16'b1001101100000100: color_data = 12'b001110100111;
		16'b1001101100000101: color_data = 12'b001110100111;
		16'b1001101100000110: color_data = 12'b001110100111;
		16'b1001101100000111: color_data = 12'b001110100111;
		16'b1001101100001000: color_data = 12'b001110100111;
		16'b1001101100001001: color_data = 12'b001110100111;
		16'b1001101100001010: color_data = 12'b001110100111;
		16'b1001101100001011: color_data = 12'b001110100111;
		16'b1001101100001100: color_data = 12'b001110100111;
		16'b1001101100001101: color_data = 12'b001110100111;
		16'b1001101100001110: color_data = 12'b001110100111;
		16'b1001101100001111: color_data = 12'b001110100111;
		16'b1001101100010000: color_data = 12'b001110100111;
		16'b1001101100010001: color_data = 12'b001110100111;
		16'b1001101100010010: color_data = 12'b001110100111;
		16'b1001101100010011: color_data = 12'b001110100111;
		16'b1001101100010100: color_data = 12'b001110100111;
		16'b1001101100010101: color_data = 12'b001110100111;
		16'b1001101100010110: color_data = 12'b001110100111;
		16'b1001101100010111: color_data = 12'b001110100111;
		16'b1001101100011000: color_data = 12'b001110100111;
		16'b1001101100011001: color_data = 12'b001110100111;
		16'b1001101100011010: color_data = 12'b001110100111;
		16'b1001101100011011: color_data = 12'b001110100111;
		16'b1001101100011100: color_data = 12'b001110100111;
		16'b1001101100011101: color_data = 12'b001110100111;
		16'b1001101100011110: color_data = 12'b001110100111;
		16'b1001101100011111: color_data = 12'b001110100111;
		16'b1001101100100000: color_data = 12'b001110100111;
		16'b1001101100100001: color_data = 12'b001110100111;
		16'b1001101100100010: color_data = 12'b001110100111;
		16'b1001101100100011: color_data = 12'b001110100111;
		16'b1001101100100100: color_data = 12'b001110100111;
		16'b1001101100100101: color_data = 12'b001110100111;
		16'b1001101100100110: color_data = 12'b001110100111;
		16'b1001101100101101: color_data = 12'b001110100111;
		16'b1001101100101110: color_data = 12'b001110100111;
		16'b1001101100101111: color_data = 12'b001110100111;
		16'b1001101100110000: color_data = 12'b001110100111;
		16'b1001101100110001: color_data = 12'b001110100111;
		16'b1001101100110010: color_data = 12'b001110100111;
		16'b1001101100110011: color_data = 12'b001110100111;
		16'b1001101100110100: color_data = 12'b001110100111;
		16'b1001101100110101: color_data = 12'b001110100111;
		16'b1001101100110110: color_data = 12'b001110100111;
		16'b1001101100110111: color_data = 12'b001110100111;
		16'b1001101100111000: color_data = 12'b001110100111;
		16'b1001101101000101: color_data = 12'b001110100111;
		16'b1001101101000110: color_data = 12'b001110100111;
		16'b1001101101000111: color_data = 12'b001110100111;
		16'b1001101101001000: color_data = 12'b001110100111;
		16'b1001101101001001: color_data = 12'b001110100111;
		16'b1001101101001010: color_data = 12'b001110100111;
		16'b1001101101001011: color_data = 12'b001110100111;
		16'b1001101101001100: color_data = 12'b001110100111;
		16'b1001101101001101: color_data = 12'b001110100111;
		16'b1001101101001110: color_data = 12'b001110100111;
		16'b1001101101001111: color_data = 12'b001110100111;
		16'b1001101101010000: color_data = 12'b001110100111;
		16'b1001101101010001: color_data = 12'b001110100111;
		16'b1001101101011000: color_data = 12'b001110100111;
		16'b1001101101011001: color_data = 12'b001110100111;
		16'b1001101101011010: color_data = 12'b001110100111;
		16'b1001101101011011: color_data = 12'b001110100111;
		16'b1001101101011100: color_data = 12'b001110100111;
		16'b1001101101011101: color_data = 12'b001110100111;
		16'b1001101101011110: color_data = 12'b001110100111;
		16'b1001101101011111: color_data = 12'b001110100111;
		16'b1001101101100000: color_data = 12'b001110100111;
		16'b1001101101100001: color_data = 12'b001110100111;
		16'b1001101101100010: color_data = 12'b001110100111;
		16'b1001101101100011: color_data = 12'b001110100111;
		16'b1001101101100100: color_data = 12'b001110100111;
		16'b1001101101100101: color_data = 12'b001110100111;
		16'b1001101101100110: color_data = 12'b001110100111;
		16'b1001101101100111: color_data = 12'b001110100111;
		16'b1001101101101000: color_data = 12'b001110100111;
		16'b1001101101101001: color_data = 12'b001110100111;
		16'b1001101101101010: color_data = 12'b001110100111;
		16'b1001101101101011: color_data = 12'b001110100111;
		16'b1001101101101100: color_data = 12'b001110100111;
		16'b1001101101101101: color_data = 12'b001110100111;
		16'b1001101101101110: color_data = 12'b001110100111;
		16'b1001101101101111: color_data = 12'b001110100111;
		16'b1001101101110000: color_data = 12'b001110100111;
		16'b1001101101110001: color_data = 12'b001110100111;
		16'b1001101101110010: color_data = 12'b001110100111;
		16'b1001101101110011: color_data = 12'b001110100111;
		16'b1001101101110100: color_data = 12'b001110100111;
		16'b1001101101110101: color_data = 12'b001110100111;
		16'b1001101101110110: color_data = 12'b001110100111;
		16'b1001101101110111: color_data = 12'b001110100111;
		16'b1001101101111000: color_data = 12'b001110100111;
		16'b1001101101111001: color_data = 12'b001110100111;
		16'b1001101101111010: color_data = 12'b001110100111;
		16'b1001101101111011: color_data = 12'b001110100111;
		16'b1001110000000000: color_data = 12'b001110100111;
		16'b1001110000000001: color_data = 12'b001110100111;
		16'b1001110000000010: color_data = 12'b001110100111;
		16'b1001110000000011: color_data = 12'b001110100111;
		16'b1001110000000100: color_data = 12'b001110100111;
		16'b1001110000000101: color_data = 12'b001110100111;
		16'b1001110000000110: color_data = 12'b001110100111;
		16'b1001110000000111: color_data = 12'b001110100111;
		16'b1001110000001000: color_data = 12'b001110100111;
		16'b1001110000001001: color_data = 12'b001110100111;
		16'b1001110000001010: color_data = 12'b001110100111;
		16'b1001110000001011: color_data = 12'b001110100111;
		16'b1001110000001100: color_data = 12'b001110100111;
		16'b1001110000001101: color_data = 12'b001110100111;
		16'b1001110000001110: color_data = 12'b001110100111;
		16'b1001110000001111: color_data = 12'b001110100111;
		16'b1001110000010000: color_data = 12'b001110100111;
		16'b1001110000010001: color_data = 12'b001110100111;
		16'b1001110000010010: color_data = 12'b001110100111;
		16'b1001110000010011: color_data = 12'b001110100111;
		16'b1001110000010100: color_data = 12'b001110100111;
		16'b1001110000010101: color_data = 12'b001110100111;
		16'b1001110000010110: color_data = 12'b001110100111;
		16'b1001110000010111: color_data = 12'b001110100111;
		16'b1001110000011000: color_data = 12'b001110100111;
		16'b1001110000011001: color_data = 12'b001110100111;
		16'b1001110000011010: color_data = 12'b001110100111;
		16'b1001110000011011: color_data = 12'b001110100111;
		16'b1001110000011100: color_data = 12'b001110100111;
		16'b1001110000011101: color_data = 12'b001110100111;
		16'b1001110000011110: color_data = 12'b001110100111;
		16'b1001110000011111: color_data = 12'b001110100111;
		16'b1001110000100000: color_data = 12'b001110100111;
		16'b1001110000100001: color_data = 12'b001110100111;
		16'b1001110000100010: color_data = 12'b001110100111;
		16'b1001110000100011: color_data = 12'b001110100111;
		16'b1001110000100100: color_data = 12'b001110100111;
		16'b1001110000101011: color_data = 12'b001110100111;
		16'b1001110000101100: color_data = 12'b001110100111;
		16'b1001110000101101: color_data = 12'b001110100111;
		16'b1001110000101110: color_data = 12'b001110100111;
		16'b1001110000101111: color_data = 12'b001110100111;
		16'b1001110000110000: color_data = 12'b001110100111;
		16'b1001110000110001: color_data = 12'b001110100111;
		16'b1001110000110010: color_data = 12'b001110100111;
		16'b1001110000110011: color_data = 12'b001110100111;
		16'b1001110000110100: color_data = 12'b001110100111;
		16'b1001110000110101: color_data = 12'b001110100111;
		16'b1001110000110110: color_data = 12'b001110100111;
		16'b1001110000110111: color_data = 12'b001110100111;
		16'b1001110001000100: color_data = 12'b001110100111;
		16'b1001110001000101: color_data = 12'b001110100111;
		16'b1001110001000110: color_data = 12'b001110100111;
		16'b1001110001000111: color_data = 12'b001110100111;
		16'b1001110001001000: color_data = 12'b001110100111;
		16'b1001110001001001: color_data = 12'b001110100111;
		16'b1001110001001010: color_data = 12'b001110100111;
		16'b1001110001001011: color_data = 12'b001110100111;
		16'b1001110001001100: color_data = 12'b001110100111;
		16'b1001110001001101: color_data = 12'b001110100111;
		16'b1001110001001110: color_data = 12'b001110100111;
		16'b1001110001001111: color_data = 12'b001110100111;
		16'b1001110001010110: color_data = 12'b001110100111;
		16'b1001110001010111: color_data = 12'b001110100111;
		16'b1001110001011000: color_data = 12'b001110100111;
		16'b1001110001011001: color_data = 12'b001110100111;
		16'b1001110001011010: color_data = 12'b001110100111;
		16'b1001110001011011: color_data = 12'b001110100111;
		16'b1001110001011100: color_data = 12'b001110100111;
		16'b1001110001011101: color_data = 12'b001110100111;
		16'b1001110001011110: color_data = 12'b001110100111;
		16'b1001110001011111: color_data = 12'b001110100111;
		16'b1001110001100000: color_data = 12'b001110100111;
		16'b1001110001100001: color_data = 12'b001110100111;
		16'b1001110001100010: color_data = 12'b001110100111;
		16'b1001110001100011: color_data = 12'b001110100111;
		16'b1001110001100100: color_data = 12'b001110100111;
		16'b1001110001100101: color_data = 12'b001110100111;
		16'b1001110001100110: color_data = 12'b001110100111;
		16'b1001110001100111: color_data = 12'b001110100111;
		16'b1001110001101000: color_data = 12'b001110100111;
		16'b1001110001101001: color_data = 12'b001110100111;
		16'b1001110001101010: color_data = 12'b001110100111;
		16'b1001110001101011: color_data = 12'b001110100111;
		16'b1001110001101100: color_data = 12'b001110100111;
		16'b1001110001101101: color_data = 12'b001110100111;
		16'b1001110001101110: color_data = 12'b001110100111;
		16'b1001110001110101: color_data = 12'b001110100111;
		16'b1001110001110110: color_data = 12'b001110100111;
		16'b1001110001110111: color_data = 12'b001110100111;
		16'b1001110001111000: color_data = 12'b001110100111;
		16'b1001110001111001: color_data = 12'b001110100111;
		16'b1001110001111010: color_data = 12'b001110100111;
		16'b1001110001111011: color_data = 12'b001110100111;
		16'b1001110001111100: color_data = 12'b001110100111;
		16'b1001110001111101: color_data = 12'b001110100111;
		16'b1001110001111110: color_data = 12'b001110100111;
		16'b1001110001111111: color_data = 12'b001110100111;
		16'b1001110010000000: color_data = 12'b001110100111;
		16'b1001110010001101: color_data = 12'b001110100111;
		16'b1001110010001110: color_data = 12'b001110100111;
		16'b1001110010001111: color_data = 12'b001110100111;
		16'b1001110010010000: color_data = 12'b001110100111;
		16'b1001110010010001: color_data = 12'b001110100111;
		16'b1001110010010010: color_data = 12'b001110100111;
		16'b1001110010010011: color_data = 12'b001110100111;
		16'b1001110010010100: color_data = 12'b001110100111;
		16'b1001110010010101: color_data = 12'b001110100111;
		16'b1001110010010110: color_data = 12'b001110100111;
		16'b1001110010010111: color_data = 12'b001110100111;
		16'b1001110010011000: color_data = 12'b001110100111;
		16'b1001110010011001: color_data = 12'b001110100111;
		16'b1001110010100000: color_data = 12'b001110100111;
		16'b1001110010100001: color_data = 12'b001110100111;
		16'b1001110010100010: color_data = 12'b001110100111;
		16'b1001110010100011: color_data = 12'b001110100111;
		16'b1001110010100100: color_data = 12'b001110100111;
		16'b1001110010100101: color_data = 12'b001110100111;
		16'b1001110010100110: color_data = 12'b001110100111;
		16'b1001110010100111: color_data = 12'b001110100111;
		16'b1001110010101000: color_data = 12'b001110100111;
		16'b1001110010101001: color_data = 12'b001110100111;
		16'b1001110010101010: color_data = 12'b001110100111;
		16'b1001110010101011: color_data = 12'b001110100111;
		16'b1001110010101100: color_data = 12'b001110100111;
		16'b1001110010101101: color_data = 12'b001110100111;
		16'b1001110010101110: color_data = 12'b001110100111;
		16'b1001110010101111: color_data = 12'b001110100111;
		16'b1001110010110000: color_data = 12'b001110100111;
		16'b1001110010110001: color_data = 12'b001110100111;
		16'b1001110010110010: color_data = 12'b001110100111;
		16'b1001110010110011: color_data = 12'b001110100111;
		16'b1001110010110100: color_data = 12'b001110100111;
		16'b1001110010110101: color_data = 12'b001110100111;
		16'b1001110010110110: color_data = 12'b001110100111;
		16'b1001110010110111: color_data = 12'b001110100111;
		16'b1001110010111000: color_data = 12'b001110100111;
		16'b1001110010111001: color_data = 12'b001110100111;
		16'b1001110010111010: color_data = 12'b001110100111;
		16'b1001110010111011: color_data = 12'b001110100111;
		16'b1001110010111100: color_data = 12'b001110100111;
		16'b1001110010111101: color_data = 12'b001110100111;
		16'b1001110010111110: color_data = 12'b001110100111;
		16'b1001110010111111: color_data = 12'b001110100111;
		16'b1001110011000000: color_data = 12'b001110100111;
		16'b1001110011000001: color_data = 12'b001110100111;
		16'b1001110011000010: color_data = 12'b001110100111;
		16'b1001110011000011: color_data = 12'b001110100111;
		16'b1001110011000100: color_data = 12'b001110100111;
		16'b1001110011001011: color_data = 12'b001110100111;
		16'b1001110011001100: color_data = 12'b001110100111;
		16'b1001110011001101: color_data = 12'b001110100111;
		16'b1001110011001110: color_data = 12'b001110100111;
		16'b1001110011001111: color_data = 12'b001110100111;
		16'b1001110011010000: color_data = 12'b001110100111;
		16'b1001110011010001: color_data = 12'b001110100111;
		16'b1001110011010010: color_data = 12'b001110100111;
		16'b1001110011010011: color_data = 12'b001110100111;
		16'b1001110011010100: color_data = 12'b001110100111;
		16'b1001110011010101: color_data = 12'b001110100111;
		16'b1001110011010110: color_data = 12'b001110100111;
		16'b1001110011110110: color_data = 12'b001110100111;
		16'b1001110011110111: color_data = 12'b001110100111;
		16'b1001110011111000: color_data = 12'b001110100111;
		16'b1001110011111001: color_data = 12'b001110100111;
		16'b1001110011111010: color_data = 12'b001110100111;
		16'b1001110011111011: color_data = 12'b001110100111;
		16'b1001110011111100: color_data = 12'b001110100111;
		16'b1001110011111101: color_data = 12'b001110100111;
		16'b1001110011111110: color_data = 12'b001110100111;
		16'b1001110011111111: color_data = 12'b001110100111;
		16'b1001110100000000: color_data = 12'b001110100111;
		16'b1001110100000001: color_data = 12'b001110100111;
		16'b1001110100000010: color_data = 12'b001110100111;
		16'b1001110100000011: color_data = 12'b001110100111;
		16'b1001110100000100: color_data = 12'b001110100111;
		16'b1001110100000101: color_data = 12'b001110100111;
		16'b1001110100000110: color_data = 12'b001110100111;
		16'b1001110100000111: color_data = 12'b001110100111;
		16'b1001110100001000: color_data = 12'b001110100111;
		16'b1001110100001001: color_data = 12'b001110100111;
		16'b1001110100001010: color_data = 12'b001110100111;
		16'b1001110100001011: color_data = 12'b001110100111;
		16'b1001110100001100: color_data = 12'b001110100111;
		16'b1001110100001101: color_data = 12'b001110100111;
		16'b1001110100001110: color_data = 12'b001110100111;
		16'b1001110100001111: color_data = 12'b001110100111;
		16'b1001110100010000: color_data = 12'b001110100111;
		16'b1001110100010001: color_data = 12'b001110100111;
		16'b1001110100010010: color_data = 12'b001110100111;
		16'b1001110100010011: color_data = 12'b001110100111;
		16'b1001110100010100: color_data = 12'b001110100111;
		16'b1001110100010101: color_data = 12'b001110100111;
		16'b1001110100010110: color_data = 12'b001110100111;
		16'b1001110100010111: color_data = 12'b001110100111;
		16'b1001110100011000: color_data = 12'b001110100111;
		16'b1001110100011001: color_data = 12'b001110100111;
		16'b1001110100011010: color_data = 12'b001110100111;
		16'b1001110100011011: color_data = 12'b001110100111;
		16'b1001110100011100: color_data = 12'b001110100111;
		16'b1001110100011101: color_data = 12'b001110100111;
		16'b1001110100011110: color_data = 12'b001110100111;
		16'b1001110100011111: color_data = 12'b001110100111;
		16'b1001110100100000: color_data = 12'b001110100111;
		16'b1001110100100001: color_data = 12'b001110100111;
		16'b1001110100100010: color_data = 12'b001110100111;
		16'b1001110100100011: color_data = 12'b001110100111;
		16'b1001110100100100: color_data = 12'b001110100111;
		16'b1001110100100101: color_data = 12'b001110100111;
		16'b1001110100100110: color_data = 12'b001110100111;
		16'b1001110100101101: color_data = 12'b001110100111;
		16'b1001110100101110: color_data = 12'b001110100111;
		16'b1001110100101111: color_data = 12'b001110100111;
		16'b1001110100110000: color_data = 12'b001110100111;
		16'b1001110100110001: color_data = 12'b001110100111;
		16'b1001110100110010: color_data = 12'b001110100111;
		16'b1001110100110011: color_data = 12'b001110100111;
		16'b1001110100110100: color_data = 12'b001110100111;
		16'b1001110100110101: color_data = 12'b001110100111;
		16'b1001110100110110: color_data = 12'b001110100111;
		16'b1001110100110111: color_data = 12'b001110100111;
		16'b1001110100111000: color_data = 12'b001110100111;
		16'b1001110101000101: color_data = 12'b001110100111;
		16'b1001110101000110: color_data = 12'b001110100111;
		16'b1001110101000111: color_data = 12'b001110100111;
		16'b1001110101001000: color_data = 12'b001110100111;
		16'b1001110101001001: color_data = 12'b001110100111;
		16'b1001110101001010: color_data = 12'b001110100111;
		16'b1001110101001011: color_data = 12'b001110100111;
		16'b1001110101001100: color_data = 12'b001110100111;
		16'b1001110101001101: color_data = 12'b001110100111;
		16'b1001110101001110: color_data = 12'b001110100111;
		16'b1001110101001111: color_data = 12'b001110100111;
		16'b1001110101010000: color_data = 12'b001110100111;
		16'b1001110101010001: color_data = 12'b001110100111;
		16'b1001110101011000: color_data = 12'b001110100111;
		16'b1001110101011001: color_data = 12'b001110100111;
		16'b1001110101011010: color_data = 12'b001110100111;
		16'b1001110101011011: color_data = 12'b001110100111;
		16'b1001110101011100: color_data = 12'b001110100111;
		16'b1001110101011101: color_data = 12'b001110100111;
		16'b1001110101011110: color_data = 12'b001110100111;
		16'b1001110101011111: color_data = 12'b001110100111;
		16'b1001110101100000: color_data = 12'b001110100111;
		16'b1001110101100001: color_data = 12'b001110100111;
		16'b1001110101100010: color_data = 12'b001110100111;
		16'b1001110101100011: color_data = 12'b001110100111;
		16'b1001110101100100: color_data = 12'b001110100111;
		16'b1001110101100101: color_data = 12'b001110100111;
		16'b1001110101100110: color_data = 12'b001110100111;
		16'b1001110101100111: color_data = 12'b001110100111;
		16'b1001110101101000: color_data = 12'b001110100111;
		16'b1001110101101001: color_data = 12'b001110100111;
		16'b1001110101101010: color_data = 12'b001110100111;
		16'b1001110101101011: color_data = 12'b001110100111;
		16'b1001110101101100: color_data = 12'b001110100111;
		16'b1001110101101101: color_data = 12'b001110100111;
		16'b1001110101101110: color_data = 12'b001110100111;
		16'b1001110101101111: color_data = 12'b001110100111;
		16'b1001110101110000: color_data = 12'b001110100111;
		16'b1001110101110001: color_data = 12'b001110100111;
		16'b1001110101110010: color_data = 12'b001110100111;
		16'b1001110101110011: color_data = 12'b001110100111;
		16'b1001110101110100: color_data = 12'b001110100111;
		16'b1001110101110101: color_data = 12'b001110100111;
		16'b1001110101110110: color_data = 12'b001110100111;
		16'b1001110101110111: color_data = 12'b001110100111;
		16'b1001110101111000: color_data = 12'b001110100111;
		16'b1001110101111001: color_data = 12'b001110100111;
		16'b1001110101111010: color_data = 12'b001110100111;
		16'b1001110101111011: color_data = 12'b001110100111;
		16'b1001111000000000: color_data = 12'b001110100111;
		16'b1001111000000001: color_data = 12'b001110100111;
		16'b1001111000000010: color_data = 12'b001110100111;
		16'b1001111000000011: color_data = 12'b001110100111;
		16'b1001111000000100: color_data = 12'b001110100111;
		16'b1001111000000101: color_data = 12'b001110100111;
		16'b1001111000000110: color_data = 12'b001110100111;
		16'b1001111000000111: color_data = 12'b001110100111;
		16'b1001111000001000: color_data = 12'b001110100111;
		16'b1001111000001001: color_data = 12'b001110100111;
		16'b1001111000001010: color_data = 12'b001110100111;
		16'b1001111000001011: color_data = 12'b001110100111;
		16'b1001111000001100: color_data = 12'b001110100111;
		16'b1001111000001101: color_data = 12'b001110100111;
		16'b1001111000001110: color_data = 12'b001110100111;
		16'b1001111000001111: color_data = 12'b001110100111;
		16'b1001111000010000: color_data = 12'b001110100111;
		16'b1001111000010001: color_data = 12'b001110100111;
		16'b1001111000010010: color_data = 12'b001110100111;
		16'b1001111000010011: color_data = 12'b001110100111;
		16'b1001111000010100: color_data = 12'b001110100111;
		16'b1001111000010101: color_data = 12'b001110100111;
		16'b1001111000010110: color_data = 12'b001110100111;
		16'b1001111000010111: color_data = 12'b001110100111;
		16'b1001111000011000: color_data = 12'b001110100111;
		16'b1001111000011001: color_data = 12'b001110100111;
		16'b1001111000011010: color_data = 12'b001110100111;
		16'b1001111000011011: color_data = 12'b001110100111;
		16'b1001111000011100: color_data = 12'b001110100111;
		16'b1001111000011101: color_data = 12'b001110100111;
		16'b1001111000011110: color_data = 12'b001110100111;
		16'b1001111000011111: color_data = 12'b001110100111;
		16'b1001111000100000: color_data = 12'b001110100111;
		16'b1001111000100001: color_data = 12'b001110100111;
		16'b1001111000100010: color_data = 12'b001110100111;
		16'b1001111000100011: color_data = 12'b001110100111;
		16'b1001111000100100: color_data = 12'b001110100111;
		16'b1001111000101011: color_data = 12'b001110100111;
		16'b1001111000101100: color_data = 12'b001110100111;
		16'b1001111000101101: color_data = 12'b001110100111;
		16'b1001111000101110: color_data = 12'b001110100111;
		16'b1001111000101111: color_data = 12'b001110100111;
		16'b1001111000110000: color_data = 12'b001110100111;
		16'b1001111000110001: color_data = 12'b001110100111;
		16'b1001111000110010: color_data = 12'b001110100111;
		16'b1001111000110011: color_data = 12'b001110100111;
		16'b1001111000110100: color_data = 12'b001110100111;
		16'b1001111000110101: color_data = 12'b001110100111;
		16'b1001111000110110: color_data = 12'b001110100111;
		16'b1001111000110111: color_data = 12'b001110100111;
		16'b1001111001000100: color_data = 12'b001110100111;
		16'b1001111001000101: color_data = 12'b001110100111;
		16'b1001111001000110: color_data = 12'b001110100111;
		16'b1001111001000111: color_data = 12'b001110100111;
		16'b1001111001001000: color_data = 12'b001110100111;
		16'b1001111001001001: color_data = 12'b001110100111;
		16'b1001111001001010: color_data = 12'b001110100111;
		16'b1001111001001011: color_data = 12'b001110100111;
		16'b1001111001001100: color_data = 12'b001110100111;
		16'b1001111001001101: color_data = 12'b001110100111;
		16'b1001111001001110: color_data = 12'b001110100111;
		16'b1001111001001111: color_data = 12'b001110100111;
		16'b1001111001010110: color_data = 12'b001110100111;
		16'b1001111001010111: color_data = 12'b001110100111;
		16'b1001111001011000: color_data = 12'b001110100111;
		16'b1001111001011001: color_data = 12'b001110100111;
		16'b1001111001011010: color_data = 12'b001110100111;
		16'b1001111001011011: color_data = 12'b001110100111;
		16'b1001111001011100: color_data = 12'b001110100111;
		16'b1001111001011101: color_data = 12'b001110100111;
		16'b1001111001011110: color_data = 12'b001110100111;
		16'b1001111001011111: color_data = 12'b001110100111;
		16'b1001111001100000: color_data = 12'b001110100111;
		16'b1001111001100001: color_data = 12'b001110100111;
		16'b1001111001100010: color_data = 12'b001110100111;
		16'b1001111001100011: color_data = 12'b001110100111;
		16'b1001111001100100: color_data = 12'b001110100111;
		16'b1001111001100101: color_data = 12'b001110100111;
		16'b1001111001100110: color_data = 12'b001110100111;
		16'b1001111001100111: color_data = 12'b001110100111;
		16'b1001111001101000: color_data = 12'b001110100111;
		16'b1001111001101001: color_data = 12'b001110100111;
		16'b1001111001101010: color_data = 12'b001110100111;
		16'b1001111001101011: color_data = 12'b001110100111;
		16'b1001111001101100: color_data = 12'b001110100111;
		16'b1001111001101101: color_data = 12'b001110100111;
		16'b1001111001101110: color_data = 12'b001110100111;
		16'b1001111001110101: color_data = 12'b001110100111;
		16'b1001111001110110: color_data = 12'b001110100111;
		16'b1001111001110111: color_data = 12'b001110100111;
		16'b1001111001111000: color_data = 12'b001110100111;
		16'b1001111001111001: color_data = 12'b001110100111;
		16'b1001111001111010: color_data = 12'b001110100111;
		16'b1001111001111011: color_data = 12'b001110100111;
		16'b1001111001111100: color_data = 12'b001110100111;
		16'b1001111001111101: color_data = 12'b001110100111;
		16'b1001111001111110: color_data = 12'b001110100111;
		16'b1001111001111111: color_data = 12'b001110100111;
		16'b1001111010000000: color_data = 12'b001110100111;
		16'b1001111010001101: color_data = 12'b001110100111;
		16'b1001111010001110: color_data = 12'b001110100111;
		16'b1001111010001111: color_data = 12'b001110100111;
		16'b1001111010010000: color_data = 12'b001110100111;
		16'b1001111010010001: color_data = 12'b001110100111;
		16'b1001111010010010: color_data = 12'b001110100111;
		16'b1001111010010011: color_data = 12'b001110100111;
		16'b1001111010010100: color_data = 12'b001110100111;
		16'b1001111010010101: color_data = 12'b001110100111;
		16'b1001111010010110: color_data = 12'b001110100111;
		16'b1001111010010111: color_data = 12'b001110100111;
		16'b1001111010011000: color_data = 12'b001110100111;
		16'b1001111010011001: color_data = 12'b001110100111;
		16'b1001111010100000: color_data = 12'b001110100111;
		16'b1001111010100001: color_data = 12'b001110100111;
		16'b1001111010100010: color_data = 12'b001110100111;
		16'b1001111010100011: color_data = 12'b001110100111;
		16'b1001111010100100: color_data = 12'b001110100111;
		16'b1001111010100101: color_data = 12'b001110100111;
		16'b1001111010100110: color_data = 12'b001110100111;
		16'b1001111010100111: color_data = 12'b001110100111;
		16'b1001111010101000: color_data = 12'b001110100111;
		16'b1001111010101001: color_data = 12'b001110100111;
		16'b1001111010101010: color_data = 12'b001110100111;
		16'b1001111010101011: color_data = 12'b001110100111;
		16'b1001111010101100: color_data = 12'b001110100111;
		16'b1001111010101101: color_data = 12'b001110100111;
		16'b1001111010101110: color_data = 12'b001110100111;
		16'b1001111010101111: color_data = 12'b001110100111;
		16'b1001111010110000: color_data = 12'b001110100111;
		16'b1001111010110001: color_data = 12'b001110100111;
		16'b1001111010110010: color_data = 12'b001110100111;
		16'b1001111010110011: color_data = 12'b001110100111;
		16'b1001111010110100: color_data = 12'b001110100111;
		16'b1001111010110101: color_data = 12'b001110100111;
		16'b1001111010110110: color_data = 12'b001110100111;
		16'b1001111010110111: color_data = 12'b001110100111;
		16'b1001111010111000: color_data = 12'b001110100111;
		16'b1001111010111001: color_data = 12'b001110100111;
		16'b1001111010111010: color_data = 12'b001110100111;
		16'b1001111010111011: color_data = 12'b001110100111;
		16'b1001111010111100: color_data = 12'b001110100111;
		16'b1001111010111101: color_data = 12'b001110100111;
		16'b1001111010111110: color_data = 12'b001110100111;
		16'b1001111010111111: color_data = 12'b001110100111;
		16'b1001111011000000: color_data = 12'b001110100111;
		16'b1001111011000001: color_data = 12'b001110100111;
		16'b1001111011000010: color_data = 12'b001110100111;
		16'b1001111011000011: color_data = 12'b001110100111;
		16'b1001111011000100: color_data = 12'b001110100111;
		16'b1001111011001011: color_data = 12'b001110100111;
		16'b1001111011001100: color_data = 12'b001110100111;
		16'b1001111011001101: color_data = 12'b001110100111;
		16'b1001111011001110: color_data = 12'b001110100111;
		16'b1001111011001111: color_data = 12'b001110100111;
		16'b1001111011010000: color_data = 12'b001110100111;
		16'b1001111011010001: color_data = 12'b001110100111;
		16'b1001111011010010: color_data = 12'b001110100111;
		16'b1001111011010011: color_data = 12'b001110100111;
		16'b1001111011010100: color_data = 12'b001110100111;
		16'b1001111011010101: color_data = 12'b001110100111;
		16'b1001111011010110: color_data = 12'b001110100111;
		16'b1001111011110110: color_data = 12'b001110100111;
		16'b1001111011110111: color_data = 12'b001110100111;
		16'b1001111011111000: color_data = 12'b001110100111;
		16'b1001111011111001: color_data = 12'b001110100111;
		16'b1001111011111010: color_data = 12'b001110100111;
		16'b1001111011111011: color_data = 12'b001110100111;
		16'b1001111011111100: color_data = 12'b001110100111;
		16'b1001111011111101: color_data = 12'b001110100111;
		16'b1001111011111110: color_data = 12'b001110100111;
		16'b1001111011111111: color_data = 12'b001110100111;
		16'b1001111100000000: color_data = 12'b001110100111;
		16'b1001111100000001: color_data = 12'b001110100111;
		16'b1001111100000010: color_data = 12'b001110100111;
		16'b1001111100000011: color_data = 12'b001110100111;
		16'b1001111100000100: color_data = 12'b001110100111;
		16'b1001111100000101: color_data = 12'b001110100111;
		16'b1001111100000110: color_data = 12'b001110100111;
		16'b1001111100000111: color_data = 12'b001110100111;
		16'b1001111100001000: color_data = 12'b001110100111;
		16'b1001111100001001: color_data = 12'b001110100111;
		16'b1001111100001010: color_data = 12'b001110100111;
		16'b1001111100001011: color_data = 12'b001110100111;
		16'b1001111100001100: color_data = 12'b001110100111;
		16'b1001111100001101: color_data = 12'b001110100111;
		16'b1001111100001110: color_data = 12'b001110100111;
		16'b1001111100001111: color_data = 12'b001110100111;
		16'b1001111100010000: color_data = 12'b001110100111;
		16'b1001111100010001: color_data = 12'b001110100111;
		16'b1001111100010010: color_data = 12'b001110100111;
		16'b1001111100010011: color_data = 12'b001110100111;
		16'b1001111100010100: color_data = 12'b001110100111;
		16'b1001111100010101: color_data = 12'b001110100111;
		16'b1001111100010110: color_data = 12'b001110100111;
		16'b1001111100010111: color_data = 12'b001110100111;
		16'b1001111100011000: color_data = 12'b001110100111;
		16'b1001111100011001: color_data = 12'b001110100111;
		16'b1001111100011010: color_data = 12'b001110100111;
		16'b1001111100011011: color_data = 12'b001110100111;
		16'b1001111100011100: color_data = 12'b001110100111;
		16'b1001111100011101: color_data = 12'b001110100111;
		16'b1001111100011110: color_data = 12'b001110100111;
		16'b1001111100011111: color_data = 12'b001110100111;
		16'b1001111100100000: color_data = 12'b001110100111;
		16'b1001111100100001: color_data = 12'b001110100111;
		16'b1001111100100010: color_data = 12'b001110100111;
		16'b1001111100100011: color_data = 12'b001110100111;
		16'b1001111100100100: color_data = 12'b001110100111;
		16'b1001111100100101: color_data = 12'b001110100111;
		16'b1001111100100110: color_data = 12'b001110100111;
		16'b1001111100101101: color_data = 12'b001110100111;
		16'b1001111100101110: color_data = 12'b001110100111;
		16'b1001111100101111: color_data = 12'b001110100111;
		16'b1001111100110000: color_data = 12'b001110100111;
		16'b1001111100110001: color_data = 12'b001110100111;
		16'b1001111100110010: color_data = 12'b001110100111;
		16'b1001111100110011: color_data = 12'b001110100111;
		16'b1001111100110100: color_data = 12'b001110100111;
		16'b1001111100110101: color_data = 12'b001110100111;
		16'b1001111100110110: color_data = 12'b001110100111;
		16'b1001111100110111: color_data = 12'b001110100111;
		16'b1001111100111000: color_data = 12'b001110100111;
		16'b1001111101000101: color_data = 12'b001110100111;
		16'b1001111101000110: color_data = 12'b001110100111;
		16'b1001111101000111: color_data = 12'b001110100111;
		16'b1001111101001000: color_data = 12'b001110100111;
		16'b1001111101001001: color_data = 12'b001110100111;
		16'b1001111101001010: color_data = 12'b001110100111;
		16'b1001111101001011: color_data = 12'b001110100111;
		16'b1001111101001100: color_data = 12'b001110100111;
		16'b1001111101001101: color_data = 12'b001110100111;
		16'b1001111101001110: color_data = 12'b001110100111;
		16'b1001111101001111: color_data = 12'b001110100111;
		16'b1001111101010000: color_data = 12'b001110100111;
		16'b1001111101010001: color_data = 12'b001110100111;
		16'b1001111101011000: color_data = 12'b001110100111;
		16'b1001111101011001: color_data = 12'b001110100111;
		16'b1001111101011010: color_data = 12'b001110100111;
		16'b1001111101011011: color_data = 12'b001110100111;
		16'b1001111101011100: color_data = 12'b001110100111;
		16'b1001111101011101: color_data = 12'b001110100111;
		16'b1001111101011110: color_data = 12'b001110100111;
		16'b1001111101011111: color_data = 12'b001110100111;
		16'b1001111101100000: color_data = 12'b001110100111;
		16'b1001111101100001: color_data = 12'b001110100111;
		16'b1001111101100010: color_data = 12'b001110100111;
		16'b1001111101100011: color_data = 12'b001110100111;
		16'b1001111101100100: color_data = 12'b001110100111;
		16'b1001111101100101: color_data = 12'b001110100111;
		16'b1001111101100110: color_data = 12'b001110100111;
		16'b1001111101100111: color_data = 12'b001110100111;
		16'b1001111101101000: color_data = 12'b001110100111;
		16'b1001111101101001: color_data = 12'b001110100111;
		16'b1001111101101010: color_data = 12'b001110100111;
		16'b1001111101101011: color_data = 12'b001110100111;
		16'b1001111101101100: color_data = 12'b001110100111;
		16'b1001111101101101: color_data = 12'b001110100111;
		16'b1001111101101110: color_data = 12'b001110100111;
		16'b1001111101101111: color_data = 12'b001110100111;
		16'b1001111101110000: color_data = 12'b001110100111;
		16'b1001111101110001: color_data = 12'b001110100111;
		16'b1001111101110010: color_data = 12'b001110100111;
		16'b1001111101110011: color_data = 12'b001110100111;
		16'b1001111101110100: color_data = 12'b001110100111;
		16'b1001111101110101: color_data = 12'b001110100111;
		16'b1001111101110110: color_data = 12'b001110100111;
		16'b1001111101110111: color_data = 12'b001110100111;
		16'b1001111101111000: color_data = 12'b001110100111;
		16'b1001111101111001: color_data = 12'b001110100111;
		16'b1001111101111010: color_data = 12'b001110100111;
		16'b1001111101111011: color_data = 12'b001110100111;
		16'b1010000000000000: color_data = 12'b001110100111;
		16'b1010000000000001: color_data = 12'b001110100111;
		16'b1010000000000010: color_data = 12'b001110100111;
		16'b1010000000000011: color_data = 12'b001110100111;
		16'b1010000000000100: color_data = 12'b001110100111;
		16'b1010000000000101: color_data = 12'b001110100111;
		16'b1010000000000110: color_data = 12'b001110100111;
		16'b1010000000000111: color_data = 12'b001110100111;
		16'b1010000000001000: color_data = 12'b001110100111;
		16'b1010000000001001: color_data = 12'b001110100111;
		16'b1010000000001010: color_data = 12'b001110100111;
		16'b1010000000001011: color_data = 12'b001110100111;
		16'b1010000000001100: color_data = 12'b001110100111;
		16'b1010000000001101: color_data = 12'b001110100111;
		16'b1010000000001110: color_data = 12'b001110100111;
		16'b1010000000001111: color_data = 12'b001110100111;
		16'b1010000000010000: color_data = 12'b001110100111;
		16'b1010000000010001: color_data = 12'b001110100111;
		16'b1010000000010010: color_data = 12'b001110100111;
		16'b1010000000010011: color_data = 12'b001110100111;
		16'b1010000000010100: color_data = 12'b001110100111;
		16'b1010000000010101: color_data = 12'b001110100111;
		16'b1010000000010110: color_data = 12'b001110100111;
		16'b1010000000010111: color_data = 12'b001110100111;
		16'b1010000000011000: color_data = 12'b001110100111;
		16'b1010000000011001: color_data = 12'b001110100111;
		16'b1010000000011010: color_data = 12'b001110100111;
		16'b1010000000011011: color_data = 12'b001110100111;
		16'b1010000000011100: color_data = 12'b001110100111;
		16'b1010000000011101: color_data = 12'b001110100111;
		16'b1010000000011110: color_data = 12'b001110100111;
		16'b1010000000011111: color_data = 12'b001110100111;
		16'b1010000000100000: color_data = 12'b001110100111;
		16'b1010000000100001: color_data = 12'b001110100111;
		16'b1010000000100010: color_data = 12'b001110100111;
		16'b1010000000100011: color_data = 12'b001110100111;
		16'b1010000000100100: color_data = 12'b001110100111;
		16'b1010000000101011: color_data = 12'b001110100111;
		16'b1010000000101100: color_data = 12'b001110100111;
		16'b1010000000101101: color_data = 12'b001110100111;
		16'b1010000000101110: color_data = 12'b001110100111;
		16'b1010000000101111: color_data = 12'b001110100111;
		16'b1010000000110000: color_data = 12'b001110100111;
		16'b1010000000110001: color_data = 12'b001110100111;
		16'b1010000000110010: color_data = 12'b001110100111;
		16'b1010000000110011: color_data = 12'b001110100111;
		16'b1010000000110100: color_data = 12'b001110100111;
		16'b1010000000110101: color_data = 12'b001110100111;
		16'b1010000000110110: color_data = 12'b001110100111;
		16'b1010000000110111: color_data = 12'b001110100111;
		16'b1010000001000100: color_data = 12'b001110100111;
		16'b1010000001000101: color_data = 12'b001110100111;
		16'b1010000001000110: color_data = 12'b001110100111;
		16'b1010000001000111: color_data = 12'b001110100111;
		16'b1010000001001000: color_data = 12'b001110100111;
		16'b1010000001001001: color_data = 12'b001110100111;
		16'b1010000001001010: color_data = 12'b001110100111;
		16'b1010000001001011: color_data = 12'b001110100111;
		16'b1010000001001100: color_data = 12'b001110100111;
		16'b1010000001001101: color_data = 12'b001110100111;
		16'b1010000001001110: color_data = 12'b001110100111;
		16'b1010000001001111: color_data = 12'b001110100111;
		16'b1010000001010110: color_data = 12'b001110100111;
		16'b1010000001010111: color_data = 12'b001110100111;
		16'b1010000001011000: color_data = 12'b001110100111;
		16'b1010000001011001: color_data = 12'b001110100111;
		16'b1010000001011010: color_data = 12'b001110100111;
		16'b1010000001011011: color_data = 12'b001110100111;
		16'b1010000001011100: color_data = 12'b001110100111;
		16'b1010000001011101: color_data = 12'b001110100111;
		16'b1010000001011110: color_data = 12'b001110100111;
		16'b1010000001011111: color_data = 12'b001110100111;
		16'b1010000001100000: color_data = 12'b001110100111;
		16'b1010000001100001: color_data = 12'b001110100111;
		16'b1010000001100010: color_data = 12'b001110100111;
		16'b1010000001100011: color_data = 12'b001110100111;
		16'b1010000001100100: color_data = 12'b001110100111;
		16'b1010000001100101: color_data = 12'b001110100111;
		16'b1010000001100110: color_data = 12'b001110100111;
		16'b1010000001100111: color_data = 12'b001110100111;
		16'b1010000001101000: color_data = 12'b001110100111;
		16'b1010000001101001: color_data = 12'b001110100111;
		16'b1010000001101010: color_data = 12'b001110100111;
		16'b1010000001101011: color_data = 12'b001110100111;
		16'b1010000001101100: color_data = 12'b001110100111;
		16'b1010000001101101: color_data = 12'b001110100111;
		16'b1010000001101110: color_data = 12'b001110100111;
		16'b1010000001110101: color_data = 12'b001110100111;
		16'b1010000001110110: color_data = 12'b001110100111;
		16'b1010000001110111: color_data = 12'b001110100111;
		16'b1010000001111000: color_data = 12'b001110100111;
		16'b1010000001111001: color_data = 12'b001110100111;
		16'b1010000001111010: color_data = 12'b001110100111;
		16'b1010000001111011: color_data = 12'b001110100111;
		16'b1010000001111100: color_data = 12'b001110100111;
		16'b1010000001111101: color_data = 12'b001110100111;
		16'b1010000001111110: color_data = 12'b001110100111;
		16'b1010000001111111: color_data = 12'b001110100111;
		16'b1010000010000000: color_data = 12'b001110100111;
		16'b1010000010001101: color_data = 12'b001110100111;
		16'b1010000010001110: color_data = 12'b001110100111;
		16'b1010000010001111: color_data = 12'b001110100111;
		16'b1010000010010000: color_data = 12'b001110100111;
		16'b1010000010010001: color_data = 12'b001110100111;
		16'b1010000010010010: color_data = 12'b001110100111;
		16'b1010000010010011: color_data = 12'b001110100111;
		16'b1010000010010100: color_data = 12'b001110100111;
		16'b1010000010010101: color_data = 12'b001110100111;
		16'b1010000010010110: color_data = 12'b001110100111;
		16'b1010000010010111: color_data = 12'b001110100111;
		16'b1010000010011000: color_data = 12'b001110100111;
		16'b1010000010011001: color_data = 12'b001110100111;
		16'b1010000010100000: color_data = 12'b001110100111;
		16'b1010000010100001: color_data = 12'b001110100111;
		16'b1010000010100010: color_data = 12'b001110100111;
		16'b1010000010100011: color_data = 12'b001110100111;
		16'b1010000010100100: color_data = 12'b001110100111;
		16'b1010000010100101: color_data = 12'b001110100111;
		16'b1010000010100110: color_data = 12'b001110100111;
		16'b1010000010100111: color_data = 12'b001110100111;
		16'b1010000010101000: color_data = 12'b001110100111;
		16'b1010000010101001: color_data = 12'b001110100111;
		16'b1010000010101010: color_data = 12'b001110100111;
		16'b1010000010101011: color_data = 12'b001110100111;
		16'b1010000010101100: color_data = 12'b001110100111;
		16'b1010000010101101: color_data = 12'b001110100111;
		16'b1010000010101110: color_data = 12'b001110100111;
		16'b1010000010101111: color_data = 12'b001110100111;
		16'b1010000010110000: color_data = 12'b001110100111;
		16'b1010000010110001: color_data = 12'b001110100111;
		16'b1010000010110010: color_data = 12'b001110100111;
		16'b1010000010110011: color_data = 12'b001110100111;
		16'b1010000010110100: color_data = 12'b001110100111;
		16'b1010000010110101: color_data = 12'b001110100111;
		16'b1010000010110110: color_data = 12'b001110100111;
		16'b1010000010110111: color_data = 12'b001110100111;
		16'b1010000010111000: color_data = 12'b001110100111;
		16'b1010000010111001: color_data = 12'b001110100111;
		16'b1010000010111010: color_data = 12'b001110100111;
		16'b1010000010111011: color_data = 12'b001110100111;
		16'b1010000010111100: color_data = 12'b001110100111;
		16'b1010000010111101: color_data = 12'b001110100111;
		16'b1010000010111110: color_data = 12'b001110100111;
		16'b1010000010111111: color_data = 12'b001110100111;
		16'b1010000011000000: color_data = 12'b001110100111;
		16'b1010000011000001: color_data = 12'b001110100111;
		16'b1010000011000010: color_data = 12'b001110100111;
		16'b1010000011000011: color_data = 12'b001110100111;
		16'b1010000011000100: color_data = 12'b001110100111;
		16'b1010000011001011: color_data = 12'b001110100111;
		16'b1010000011001100: color_data = 12'b001110100111;
		16'b1010000011001101: color_data = 12'b001110100111;
		16'b1010000011001110: color_data = 12'b001110100111;
		16'b1010000011001111: color_data = 12'b001110100111;
		16'b1010000011010000: color_data = 12'b001110100111;
		16'b1010000011010001: color_data = 12'b001110100111;
		16'b1010000011010010: color_data = 12'b001110100111;
		16'b1010000011010011: color_data = 12'b001110100111;
		16'b1010000011010100: color_data = 12'b001110100111;
		16'b1010000011010101: color_data = 12'b001110100111;
		16'b1010000011010110: color_data = 12'b001110100111;
		16'b1010000011110110: color_data = 12'b001110100111;
		16'b1010000011110111: color_data = 12'b001110100111;
		16'b1010000011111000: color_data = 12'b001110100111;
		16'b1010000011111001: color_data = 12'b001110100111;
		16'b1010000011111010: color_data = 12'b001110100111;
		16'b1010000011111011: color_data = 12'b001110100111;
		16'b1010000011111100: color_data = 12'b001110100111;
		16'b1010000011111101: color_data = 12'b001110100111;
		16'b1010000011111110: color_data = 12'b001110100111;
		16'b1010000011111111: color_data = 12'b001110100111;
		16'b1010000100000000: color_data = 12'b001110100111;
		16'b1010000100000001: color_data = 12'b001110100111;
		16'b1010000100000010: color_data = 12'b001110100111;
		16'b1010000100000011: color_data = 12'b001110100111;
		16'b1010000100000100: color_data = 12'b001110100111;
		16'b1010000100000101: color_data = 12'b001110100111;
		16'b1010000100000110: color_data = 12'b001110100111;
		16'b1010000100000111: color_data = 12'b001110100111;
		16'b1010000100001000: color_data = 12'b001110100111;
		16'b1010000100001001: color_data = 12'b001110100111;
		16'b1010000100001010: color_data = 12'b001110100111;
		16'b1010000100001011: color_data = 12'b001110100111;
		16'b1010000100001100: color_data = 12'b001110100111;
		16'b1010000100001101: color_data = 12'b001110100111;
		16'b1010000100001110: color_data = 12'b001110100111;
		16'b1010000100001111: color_data = 12'b001110100111;
		16'b1010000100010000: color_data = 12'b001110100111;
		16'b1010000100010001: color_data = 12'b001110100111;
		16'b1010000100010010: color_data = 12'b001110100111;
		16'b1010000100010011: color_data = 12'b001110100111;
		16'b1010000100010100: color_data = 12'b001110100111;
		16'b1010000100010101: color_data = 12'b001110100111;
		16'b1010000100010110: color_data = 12'b001110100111;
		16'b1010000100010111: color_data = 12'b001110100111;
		16'b1010000100011000: color_data = 12'b001110100111;
		16'b1010000100011001: color_data = 12'b001110100111;
		16'b1010000100011010: color_data = 12'b001110100111;
		16'b1010000100011011: color_data = 12'b001110100111;
		16'b1010000100011100: color_data = 12'b001110100111;
		16'b1010000100011101: color_data = 12'b001110100111;
		16'b1010000100011110: color_data = 12'b001110100111;
		16'b1010000100011111: color_data = 12'b001110100111;
		16'b1010000100100000: color_data = 12'b001110100111;
		16'b1010000100100001: color_data = 12'b001110100111;
		16'b1010000100100010: color_data = 12'b001110100111;
		16'b1010000100100011: color_data = 12'b001110100111;
		16'b1010000100100100: color_data = 12'b001110100111;
		16'b1010000100100101: color_data = 12'b001110100111;
		16'b1010000100100110: color_data = 12'b001110100111;
		16'b1010000100101101: color_data = 12'b001110100111;
		16'b1010000100101110: color_data = 12'b001110100111;
		16'b1010000100101111: color_data = 12'b001110100111;
		16'b1010000100110000: color_data = 12'b001110100111;
		16'b1010000100110001: color_data = 12'b001110100111;
		16'b1010000100110010: color_data = 12'b001110100111;
		16'b1010000100110011: color_data = 12'b001110100111;
		16'b1010000100110100: color_data = 12'b001110100111;
		16'b1010000100110101: color_data = 12'b001110100111;
		16'b1010000100110110: color_data = 12'b001110100111;
		16'b1010000100110111: color_data = 12'b001110100111;
		16'b1010000100111000: color_data = 12'b001110100111;
		16'b1010000101000101: color_data = 12'b001110100111;
		16'b1010000101000110: color_data = 12'b001110100111;
		16'b1010000101000111: color_data = 12'b001110100111;
		16'b1010000101001000: color_data = 12'b001110100111;
		16'b1010000101001001: color_data = 12'b001110100111;
		16'b1010000101001010: color_data = 12'b001110100111;
		16'b1010000101001011: color_data = 12'b001110100111;
		16'b1010000101001100: color_data = 12'b001110100111;
		16'b1010000101001101: color_data = 12'b001110100111;
		16'b1010000101001110: color_data = 12'b001110100111;
		16'b1010000101001111: color_data = 12'b001110100111;
		16'b1010000101010000: color_data = 12'b001110100111;
		16'b1010000101010001: color_data = 12'b001110100111;
		16'b1010000101011000: color_data = 12'b001110100111;
		16'b1010000101011001: color_data = 12'b001110100111;
		16'b1010000101011010: color_data = 12'b001110100111;
		16'b1010000101011011: color_data = 12'b001110100111;
		16'b1010000101011100: color_data = 12'b001110100111;
		16'b1010000101011101: color_data = 12'b001110100111;
		16'b1010000101011110: color_data = 12'b001110100111;
		16'b1010000101011111: color_data = 12'b001110100111;
		16'b1010000101100000: color_data = 12'b001110100111;
		16'b1010000101100001: color_data = 12'b001110100111;
		16'b1010000101100010: color_data = 12'b001110100111;
		16'b1010000101100011: color_data = 12'b001110100111;
		16'b1010000101100100: color_data = 12'b001110100111;
		16'b1010000101100101: color_data = 12'b001110100111;
		16'b1010000101100110: color_data = 12'b001110100111;
		16'b1010000101100111: color_data = 12'b001110100111;
		16'b1010000101101000: color_data = 12'b001110100111;
		16'b1010000101101001: color_data = 12'b001110100111;
		16'b1010000101101010: color_data = 12'b001110100111;
		16'b1010000101101011: color_data = 12'b001110100111;
		16'b1010000101101100: color_data = 12'b001110100111;
		16'b1010000101101101: color_data = 12'b001110100111;
		16'b1010000101101110: color_data = 12'b001110100111;
		16'b1010000101101111: color_data = 12'b001110100111;
		16'b1010000101110000: color_data = 12'b001110100111;
		16'b1010000101110001: color_data = 12'b001110100111;
		16'b1010000101110010: color_data = 12'b001110100111;
		16'b1010000101110011: color_data = 12'b001110100111;
		16'b1010000101110100: color_data = 12'b001110100111;
		16'b1010000101110101: color_data = 12'b001110100111;
		16'b1010000101110110: color_data = 12'b001110100111;
		16'b1010000101110111: color_data = 12'b001110100111;
		16'b1010000101111000: color_data = 12'b001110100111;
		16'b1010000101111001: color_data = 12'b001110100111;
		16'b1010000101111010: color_data = 12'b001110100111;
		16'b1010000101111011: color_data = 12'b001110100111;
		16'b1010001000000000: color_data = 12'b001110100111;
		16'b1010001000000001: color_data = 12'b001110100111;
		16'b1010001000000010: color_data = 12'b001110100111;
		16'b1010001000000011: color_data = 12'b001110100111;
		16'b1010001000000100: color_data = 12'b001110100111;
		16'b1010001000000101: color_data = 12'b001110100111;
		16'b1010001000000110: color_data = 12'b001110100111;
		16'b1010001000000111: color_data = 12'b001110100111;
		16'b1010001000001000: color_data = 12'b001110100111;
		16'b1010001000001001: color_data = 12'b001110100111;
		16'b1010001000001010: color_data = 12'b001110100111;
		16'b1010001000001011: color_data = 12'b001110100111;
		16'b1010001000001100: color_data = 12'b001110100111;
		16'b1010001000001101: color_data = 12'b001110100111;
		16'b1010001000001110: color_data = 12'b001110100111;
		16'b1010001000001111: color_data = 12'b001110100111;
		16'b1010001000010000: color_data = 12'b001110100111;
		16'b1010001000010001: color_data = 12'b001110100111;
		16'b1010001000010010: color_data = 12'b001110100111;
		16'b1010001000010011: color_data = 12'b001110100111;
		16'b1010001000010100: color_data = 12'b001110100111;
		16'b1010001000010101: color_data = 12'b001110100111;
		16'b1010001000010110: color_data = 12'b001110100111;
		16'b1010001000010111: color_data = 12'b001110100111;
		16'b1010001000011000: color_data = 12'b001110100111;
		16'b1010001000011001: color_data = 12'b001110100111;
		16'b1010001000011010: color_data = 12'b001110100111;
		16'b1010001000011011: color_data = 12'b001110100111;
		16'b1010001000011100: color_data = 12'b001110100111;
		16'b1010001000011101: color_data = 12'b001110100111;
		16'b1010001000011110: color_data = 12'b001110100111;
		16'b1010001000011111: color_data = 12'b001110100111;
		16'b1010001000100000: color_data = 12'b001110100111;
		16'b1010001000100001: color_data = 12'b001110100111;
		16'b1010001000100010: color_data = 12'b001110100111;
		16'b1010001000100011: color_data = 12'b001110100111;
		16'b1010001000100100: color_data = 12'b001110100111;
		16'b1010001000101011: color_data = 12'b001110100111;
		16'b1010001000101100: color_data = 12'b001110100111;
		16'b1010001000101101: color_data = 12'b001110100111;
		16'b1010001000101110: color_data = 12'b001110100111;
		16'b1010001000101111: color_data = 12'b001110100111;
		16'b1010001000110000: color_data = 12'b001110100111;
		16'b1010001000110001: color_data = 12'b001110100111;
		16'b1010001000110010: color_data = 12'b001110100111;
		16'b1010001000110011: color_data = 12'b001110100111;
		16'b1010001000110100: color_data = 12'b001110100111;
		16'b1010001000110101: color_data = 12'b001110100111;
		16'b1010001000110110: color_data = 12'b001110100111;
		16'b1010001000110111: color_data = 12'b001110100111;
		16'b1010001001000100: color_data = 12'b001110100111;
		16'b1010001001000101: color_data = 12'b001110100111;
		16'b1010001001000110: color_data = 12'b001110100111;
		16'b1010001001000111: color_data = 12'b001110100111;
		16'b1010001001001000: color_data = 12'b001110100111;
		16'b1010001001001001: color_data = 12'b001110100111;
		16'b1010001001001010: color_data = 12'b001110100111;
		16'b1010001001001011: color_data = 12'b001110100111;
		16'b1010001001001100: color_data = 12'b001110100111;
		16'b1010001001001101: color_data = 12'b001110100111;
		16'b1010001001001110: color_data = 12'b001110100111;
		16'b1010001001001111: color_data = 12'b001110100111;
		16'b1010001001010110: color_data = 12'b001110100111;
		16'b1010001001010111: color_data = 12'b001110100111;
		16'b1010001001011000: color_data = 12'b001110100111;
		16'b1010001001011001: color_data = 12'b001110100111;
		16'b1010001001011010: color_data = 12'b001110100111;
		16'b1010001001011011: color_data = 12'b001110100111;
		16'b1010001001011100: color_data = 12'b001110100111;
		16'b1010001001011101: color_data = 12'b001110100111;
		16'b1010001001011110: color_data = 12'b001110100111;
		16'b1010001001011111: color_data = 12'b001110100111;
		16'b1010001001100000: color_data = 12'b001110100111;
		16'b1010001001100001: color_data = 12'b001110100111;
		16'b1010001001100010: color_data = 12'b001110100111;
		16'b1010001001100011: color_data = 12'b001110100111;
		16'b1010001001100100: color_data = 12'b001110100111;
		16'b1010001001100101: color_data = 12'b001110100111;
		16'b1010001001100110: color_data = 12'b001110100111;
		16'b1010001001100111: color_data = 12'b001110100111;
		16'b1010001001101000: color_data = 12'b001110100111;
		16'b1010001001101001: color_data = 12'b001110100111;
		16'b1010001001101010: color_data = 12'b001110100111;
		16'b1010001001101011: color_data = 12'b001110100111;
		16'b1010001001101100: color_data = 12'b001110100111;
		16'b1010001001101101: color_data = 12'b001110100111;
		16'b1010001001101110: color_data = 12'b001110100111;
		16'b1010001001110101: color_data = 12'b001110100111;
		16'b1010001001110110: color_data = 12'b001110100111;
		16'b1010001001110111: color_data = 12'b001110100111;
		16'b1010001001111000: color_data = 12'b001110100111;
		16'b1010001001111001: color_data = 12'b001110100111;
		16'b1010001001111010: color_data = 12'b001110100111;
		16'b1010001001111011: color_data = 12'b001110100111;
		16'b1010001001111100: color_data = 12'b001110100111;
		16'b1010001001111101: color_data = 12'b001110100111;
		16'b1010001001111110: color_data = 12'b001110100111;
		16'b1010001001111111: color_data = 12'b001110100111;
		16'b1010001010000000: color_data = 12'b001110100111;
		16'b1010001010001101: color_data = 12'b001110100111;
		16'b1010001010001110: color_data = 12'b001110100111;
		16'b1010001010001111: color_data = 12'b001110100111;
		16'b1010001010010000: color_data = 12'b001110100111;
		16'b1010001010010001: color_data = 12'b001110100111;
		16'b1010001010010010: color_data = 12'b001110100111;
		16'b1010001010010011: color_data = 12'b001110100111;
		16'b1010001010010100: color_data = 12'b001110100111;
		16'b1010001010010101: color_data = 12'b001110100111;
		16'b1010001010010110: color_data = 12'b001110100111;
		16'b1010001010010111: color_data = 12'b001110100111;
		16'b1010001010011000: color_data = 12'b001110100111;
		16'b1010001010011001: color_data = 12'b001110100111;
		16'b1010001010100000: color_data = 12'b001110100111;
		16'b1010001010100001: color_data = 12'b001110100111;
		16'b1010001010100010: color_data = 12'b001110100111;
		16'b1010001010100011: color_data = 12'b001110100111;
		16'b1010001010100100: color_data = 12'b001110100111;
		16'b1010001010100101: color_data = 12'b001110100111;
		16'b1010001010100110: color_data = 12'b001110100111;
		16'b1010001010100111: color_data = 12'b001110100111;
		16'b1010001010101000: color_data = 12'b001110100111;
		16'b1010001010101001: color_data = 12'b001110100111;
		16'b1010001010101010: color_data = 12'b001110100111;
		16'b1010001010101011: color_data = 12'b001110100111;
		16'b1010001010101100: color_data = 12'b001110100111;
		16'b1010001010101101: color_data = 12'b001110100111;
		16'b1010001010101110: color_data = 12'b001110100111;
		16'b1010001010101111: color_data = 12'b001110100111;
		16'b1010001010110000: color_data = 12'b001110100111;
		16'b1010001010110001: color_data = 12'b001110100111;
		16'b1010001010110010: color_data = 12'b001110100111;
		16'b1010001010110011: color_data = 12'b001110100111;
		16'b1010001010110100: color_data = 12'b001110100111;
		16'b1010001010110101: color_data = 12'b001110100111;
		16'b1010001010110110: color_data = 12'b001110100111;
		16'b1010001010110111: color_data = 12'b001110100111;
		16'b1010001010111000: color_data = 12'b001110100111;
		16'b1010001010111001: color_data = 12'b001110100111;
		16'b1010001010111010: color_data = 12'b001110100111;
		16'b1010001010111011: color_data = 12'b001110100111;
		16'b1010001010111100: color_data = 12'b001110100111;
		16'b1010001010111101: color_data = 12'b001110100111;
		16'b1010001010111110: color_data = 12'b001110100111;
		16'b1010001010111111: color_data = 12'b001110100111;
		16'b1010001011000000: color_data = 12'b001110100111;
		16'b1010001011000001: color_data = 12'b001110100111;
		16'b1010001011000010: color_data = 12'b001110100111;
		16'b1010001011000011: color_data = 12'b001110100111;
		16'b1010001011000100: color_data = 12'b001110100111;
		16'b1010001011001011: color_data = 12'b001110100111;
		16'b1010001011001100: color_data = 12'b001110100111;
		16'b1010001011001101: color_data = 12'b001110100111;
		16'b1010001011001110: color_data = 12'b001110100111;
		16'b1010001011001111: color_data = 12'b001110100111;
		16'b1010001011010000: color_data = 12'b001110100111;
		16'b1010001011010001: color_data = 12'b001110100111;
		16'b1010001011010010: color_data = 12'b001110100111;
		16'b1010001011010011: color_data = 12'b001110100111;
		16'b1010001011010100: color_data = 12'b001110100111;
		16'b1010001011010101: color_data = 12'b001110100111;
		16'b1010001011010110: color_data = 12'b001110100111;
		16'b1010001011110110: color_data = 12'b001110100111;
		16'b1010001011110111: color_data = 12'b001110100111;
		16'b1010001011111000: color_data = 12'b001110100111;
		16'b1010001011111001: color_data = 12'b001110100111;
		16'b1010001011111010: color_data = 12'b001110100111;
		16'b1010001011111011: color_data = 12'b001110100111;
		16'b1010001011111100: color_data = 12'b001110100111;
		16'b1010001011111101: color_data = 12'b001110100111;
		16'b1010001011111110: color_data = 12'b001110100111;
		16'b1010001011111111: color_data = 12'b001110100111;
		16'b1010001100000000: color_data = 12'b001110100111;
		16'b1010001100000001: color_data = 12'b001110100111;
		16'b1010001100000010: color_data = 12'b001110100111;
		16'b1010001100000011: color_data = 12'b001110100111;
		16'b1010001100000100: color_data = 12'b001110100111;
		16'b1010001100000101: color_data = 12'b001110100111;
		16'b1010001100000110: color_data = 12'b001110100111;
		16'b1010001100000111: color_data = 12'b001110100111;
		16'b1010001100001000: color_data = 12'b001110100111;
		16'b1010001100001001: color_data = 12'b001110100111;
		16'b1010001100001010: color_data = 12'b001110100111;
		16'b1010001100001011: color_data = 12'b001110100111;
		16'b1010001100001100: color_data = 12'b001110100111;
		16'b1010001100001101: color_data = 12'b001110100111;
		16'b1010001100001110: color_data = 12'b001110100111;
		16'b1010001100001111: color_data = 12'b001110100111;
		16'b1010001100010000: color_data = 12'b001110100111;
		16'b1010001100010001: color_data = 12'b001110100111;
		16'b1010001100010010: color_data = 12'b001110100111;
		16'b1010001100010011: color_data = 12'b001110100111;
		16'b1010001100010100: color_data = 12'b001110100111;
		16'b1010001100010101: color_data = 12'b001110100111;
		16'b1010001100010110: color_data = 12'b001110100111;
		16'b1010001100010111: color_data = 12'b001110100111;
		16'b1010001100011000: color_data = 12'b001110100111;
		16'b1010001100011001: color_data = 12'b001110100111;
		16'b1010001100011010: color_data = 12'b001110100111;
		16'b1010001100011011: color_data = 12'b001110100111;
		16'b1010001100011100: color_data = 12'b001110100111;
		16'b1010001100011101: color_data = 12'b001110100111;
		16'b1010001100011110: color_data = 12'b001110100111;
		16'b1010001100011111: color_data = 12'b001110100111;
		16'b1010001100100000: color_data = 12'b001110100111;
		16'b1010001100100001: color_data = 12'b001110100111;
		16'b1010001100100010: color_data = 12'b001110100111;
		16'b1010001100100011: color_data = 12'b001110100111;
		16'b1010001100100100: color_data = 12'b001110100111;
		16'b1010001100100101: color_data = 12'b001110100111;
		16'b1010001100100110: color_data = 12'b001110100111;
		16'b1010001100101101: color_data = 12'b001110100111;
		16'b1010001100101110: color_data = 12'b001110100111;
		16'b1010001100101111: color_data = 12'b001110100111;
		16'b1010001100110000: color_data = 12'b001110100111;
		16'b1010001100110001: color_data = 12'b001110100111;
		16'b1010001100110010: color_data = 12'b001110100111;
		16'b1010001100110011: color_data = 12'b001110100111;
		16'b1010001100110100: color_data = 12'b001110100111;
		16'b1010001100110101: color_data = 12'b001110100111;
		16'b1010001100110110: color_data = 12'b001110100111;
		16'b1010001100110111: color_data = 12'b001110100111;
		16'b1010001100111000: color_data = 12'b001110100111;
		16'b1010001101000101: color_data = 12'b001110100111;
		16'b1010001101000110: color_data = 12'b001110100111;
		16'b1010001101000111: color_data = 12'b001110100111;
		16'b1010001101001000: color_data = 12'b001110100111;
		16'b1010001101001001: color_data = 12'b001110100111;
		16'b1010001101001010: color_data = 12'b001110100111;
		16'b1010001101001011: color_data = 12'b001110100111;
		16'b1010001101001100: color_data = 12'b001110100111;
		16'b1010001101001101: color_data = 12'b001110100111;
		16'b1010001101001110: color_data = 12'b001110100111;
		16'b1010001101001111: color_data = 12'b001110100111;
		16'b1010001101010000: color_data = 12'b001110100111;
		16'b1010001101010001: color_data = 12'b001110100111;
		16'b1010001101011000: color_data = 12'b001110100111;
		16'b1010001101011001: color_data = 12'b001110100111;
		16'b1010001101011010: color_data = 12'b001110100111;
		16'b1010001101011011: color_data = 12'b001110100111;
		16'b1010001101011100: color_data = 12'b001110100111;
		16'b1010001101011101: color_data = 12'b001110100111;
		16'b1010001101011110: color_data = 12'b001110100111;
		16'b1010001101011111: color_data = 12'b001110100111;
		16'b1010001101100000: color_data = 12'b001110100111;
		16'b1010001101100001: color_data = 12'b001110100111;
		16'b1010001101100010: color_data = 12'b001110100111;
		16'b1010001101100011: color_data = 12'b001110100111;
		16'b1010001101100100: color_data = 12'b001110100111;
		16'b1010001101100101: color_data = 12'b001110100111;
		16'b1010001101100110: color_data = 12'b001110100111;
		16'b1010001101100111: color_data = 12'b001110100111;
		16'b1010001101101000: color_data = 12'b001110100111;
		16'b1010001101101001: color_data = 12'b001110100111;
		16'b1010001101101010: color_data = 12'b001110100111;
		16'b1010001101101011: color_data = 12'b001110100111;
		16'b1010001101101100: color_data = 12'b001110100111;
		16'b1010001101101101: color_data = 12'b001110100111;
		16'b1010001101101110: color_data = 12'b001110100111;
		16'b1010001101101111: color_data = 12'b001110100111;
		16'b1010001101110000: color_data = 12'b001110100111;
		16'b1010001101110001: color_data = 12'b001110100111;
		16'b1010001101110010: color_data = 12'b001110100111;
		16'b1010001101110011: color_data = 12'b001110100111;
		16'b1010001101110100: color_data = 12'b001110100111;
		16'b1010001101110101: color_data = 12'b001110100111;
		16'b1010001101110110: color_data = 12'b001110100111;
		16'b1010001101110111: color_data = 12'b001110100111;
		16'b1010001101111000: color_data = 12'b001110100111;
		16'b1010001101111001: color_data = 12'b001110100111;
		16'b1010001101111010: color_data = 12'b001110100111;
		16'b1010001101111011: color_data = 12'b001110100111;
		16'b1010010000000000: color_data = 12'b001110100111;
		16'b1010010000000001: color_data = 12'b001110100111;
		16'b1010010000000010: color_data = 12'b001110100111;
		16'b1010010000000011: color_data = 12'b001110100111;
		16'b1010010000000100: color_data = 12'b001110100111;
		16'b1010010000000101: color_data = 12'b001110100111;
		16'b1010010000000110: color_data = 12'b001110100111;
		16'b1010010000000111: color_data = 12'b001110100111;
		16'b1010010000001000: color_data = 12'b001110100111;
		16'b1010010000001001: color_data = 12'b001110100111;
		16'b1010010000001010: color_data = 12'b001110100111;
		16'b1010010000001011: color_data = 12'b001110100111;
		16'b1010010000001100: color_data = 12'b001110100111;
		16'b1010010000001101: color_data = 12'b001110100111;
		16'b1010010000001110: color_data = 12'b001110100111;
		16'b1010010000001111: color_data = 12'b001110100111;
		16'b1010010000010000: color_data = 12'b001110100111;
		16'b1010010000010001: color_data = 12'b001110100111;
		16'b1010010000010010: color_data = 12'b001110100111;
		16'b1010010000010011: color_data = 12'b001110100111;
		16'b1010010000010100: color_data = 12'b001110100111;
		16'b1010010000010101: color_data = 12'b001110100111;
		16'b1010010000010110: color_data = 12'b001110100111;
		16'b1010010000010111: color_data = 12'b001110100111;
		16'b1010010000011000: color_data = 12'b001110100111;
		16'b1010010000011001: color_data = 12'b001110100111;
		16'b1010010000011010: color_data = 12'b001110100111;
		16'b1010010000011011: color_data = 12'b001110100111;
		16'b1010010000011100: color_data = 12'b001110100111;
		16'b1010010000011101: color_data = 12'b001110100111;
		16'b1010010000011110: color_data = 12'b001110100111;
		16'b1010010000011111: color_data = 12'b001110100111;
		16'b1010010000100000: color_data = 12'b001110100111;
		16'b1010010000100001: color_data = 12'b001110100111;
		16'b1010010000100010: color_data = 12'b001110100111;
		16'b1010010000100011: color_data = 12'b001110100111;
		16'b1010010000100100: color_data = 12'b001110100111;
		16'b1010010000101011: color_data = 12'b001110100111;
		16'b1010010000101100: color_data = 12'b001110100111;
		16'b1010010000101101: color_data = 12'b001110100111;
		16'b1010010000101110: color_data = 12'b001110100111;
		16'b1010010000101111: color_data = 12'b001110100111;
		16'b1010010000110000: color_data = 12'b001110100111;
		16'b1010010000110001: color_data = 12'b001110100111;
		16'b1010010000110010: color_data = 12'b001110100111;
		16'b1010010000110011: color_data = 12'b001110100111;
		16'b1010010000110100: color_data = 12'b001110100111;
		16'b1010010000110101: color_data = 12'b001110100111;
		16'b1010010000110110: color_data = 12'b001110100111;
		16'b1010010000110111: color_data = 12'b001110100111;
		16'b1010010001000100: color_data = 12'b001110100111;
		16'b1010010001000101: color_data = 12'b001110100111;
		16'b1010010001000110: color_data = 12'b001110100111;
		16'b1010010001000111: color_data = 12'b001110100111;
		16'b1010010001001000: color_data = 12'b001110100111;
		16'b1010010001001001: color_data = 12'b001110100111;
		16'b1010010001001010: color_data = 12'b001110100111;
		16'b1010010001001011: color_data = 12'b001110100111;
		16'b1010010001001100: color_data = 12'b001110100111;
		16'b1010010001001101: color_data = 12'b001110100111;
		16'b1010010001001110: color_data = 12'b001110100111;
		16'b1010010001001111: color_data = 12'b001110100111;
		16'b1010010001010110: color_data = 12'b001110100111;
		16'b1010010001010111: color_data = 12'b001110100111;
		16'b1010010001011000: color_data = 12'b001110100111;
		16'b1010010001011001: color_data = 12'b001110100111;
		16'b1010010001011010: color_data = 12'b001110100111;
		16'b1010010001011011: color_data = 12'b001110100111;
		16'b1010010001011100: color_data = 12'b001110100111;
		16'b1010010001011101: color_data = 12'b001110100111;
		16'b1010010001011110: color_data = 12'b001110100111;
		16'b1010010001011111: color_data = 12'b001110100111;
		16'b1010010001100000: color_data = 12'b001110100111;
		16'b1010010001100001: color_data = 12'b001110100111;
		16'b1010010001100010: color_data = 12'b001110100111;
		16'b1010010001100011: color_data = 12'b001110100111;
		16'b1010010001100100: color_data = 12'b001110100111;
		16'b1010010001100101: color_data = 12'b001110100111;
		16'b1010010001100110: color_data = 12'b001110100111;
		16'b1010010001100111: color_data = 12'b001110100111;
		16'b1010010001101000: color_data = 12'b001110100111;
		16'b1010010001101001: color_data = 12'b001110100111;
		16'b1010010001101010: color_data = 12'b001110100111;
		16'b1010010001101011: color_data = 12'b001110100111;
		16'b1010010001101100: color_data = 12'b001110100111;
		16'b1010010001101101: color_data = 12'b001110100111;
		16'b1010010001101110: color_data = 12'b001110100111;
		16'b1010010001110101: color_data = 12'b001110100111;
		16'b1010010001110110: color_data = 12'b001110100111;
		16'b1010010001110111: color_data = 12'b001110100111;
		16'b1010010001111000: color_data = 12'b001110100111;
		16'b1010010001111001: color_data = 12'b001110100111;
		16'b1010010001111010: color_data = 12'b001110100111;
		16'b1010010001111011: color_data = 12'b001110100111;
		16'b1010010001111100: color_data = 12'b001110100111;
		16'b1010010001111101: color_data = 12'b001110100111;
		16'b1010010001111110: color_data = 12'b001110100111;
		16'b1010010001111111: color_data = 12'b001110100111;
		16'b1010010010000000: color_data = 12'b001110100111;
		16'b1010010010001101: color_data = 12'b001110100111;
		16'b1010010010001110: color_data = 12'b001110100111;
		16'b1010010010001111: color_data = 12'b001110100111;
		16'b1010010010010000: color_data = 12'b001110100111;
		16'b1010010010010001: color_data = 12'b001110100111;
		16'b1010010010010010: color_data = 12'b001110100111;
		16'b1010010010010011: color_data = 12'b001110100111;
		16'b1010010010010100: color_data = 12'b001110100111;
		16'b1010010010010101: color_data = 12'b001110100111;
		16'b1010010010010110: color_data = 12'b001110100111;
		16'b1010010010010111: color_data = 12'b001110100111;
		16'b1010010010011000: color_data = 12'b001110100111;
		16'b1010010010011001: color_data = 12'b001110100111;
		16'b1010010010100000: color_data = 12'b001110100111;
		16'b1010010010100001: color_data = 12'b001110100111;
		16'b1010010010100010: color_data = 12'b001110100111;
		16'b1010010010100011: color_data = 12'b001110100111;
		16'b1010010010100100: color_data = 12'b001110100111;
		16'b1010010010100101: color_data = 12'b001110100111;
		16'b1010010010100110: color_data = 12'b001110100111;
		16'b1010010010100111: color_data = 12'b001110100111;
		16'b1010010010101000: color_data = 12'b001110100111;
		16'b1010010010101001: color_data = 12'b001110100111;
		16'b1010010010101010: color_data = 12'b001110100111;
		16'b1010010010101011: color_data = 12'b001110100111;
		16'b1010010010101100: color_data = 12'b001110100111;
		16'b1010010010101101: color_data = 12'b001110100111;
		16'b1010010010101110: color_data = 12'b001110100111;
		16'b1010010010101111: color_data = 12'b001110100111;
		16'b1010010010110000: color_data = 12'b001110100111;
		16'b1010010010110001: color_data = 12'b001110100111;
		16'b1010010010110010: color_data = 12'b001110100111;
		16'b1010010010110011: color_data = 12'b001110100111;
		16'b1010010010110100: color_data = 12'b001110100111;
		16'b1010010010110101: color_data = 12'b001110100111;
		16'b1010010010110110: color_data = 12'b001110100111;
		16'b1010010010110111: color_data = 12'b001110100111;
		16'b1010010010111000: color_data = 12'b001110100111;
		16'b1010010010111001: color_data = 12'b001110100111;
		16'b1010010010111010: color_data = 12'b001110100111;
		16'b1010010010111011: color_data = 12'b001110100111;
		16'b1010010010111100: color_data = 12'b001110100111;
		16'b1010010010111101: color_data = 12'b001110100111;
		16'b1010010010111110: color_data = 12'b001110100111;
		16'b1010010010111111: color_data = 12'b001110100111;
		16'b1010010011000000: color_data = 12'b001110100111;
		16'b1010010011000001: color_data = 12'b001110100111;
		16'b1010010011000010: color_data = 12'b001110100111;
		16'b1010010011000011: color_data = 12'b001110100111;
		16'b1010010011000100: color_data = 12'b001110100111;
		16'b1010010011001011: color_data = 12'b001110100111;
		16'b1010010011001100: color_data = 12'b001110100111;
		16'b1010010011001101: color_data = 12'b001110100111;
		16'b1010010011001110: color_data = 12'b001110100111;
		16'b1010010011001111: color_data = 12'b001110100111;
		16'b1010010011010000: color_data = 12'b001110100111;
		16'b1010010011010001: color_data = 12'b001110100111;
		16'b1010010011010010: color_data = 12'b001110100111;
		16'b1010010011010011: color_data = 12'b001110100111;
		16'b1010010011010100: color_data = 12'b001110100111;
		16'b1010010011010101: color_data = 12'b001110100111;
		16'b1010010011010110: color_data = 12'b001110100111;
		16'b1010010011110110: color_data = 12'b001110100111;
		16'b1010010011110111: color_data = 12'b001110100111;
		16'b1010010011111000: color_data = 12'b001110100111;
		16'b1010010011111001: color_data = 12'b001110100111;
		16'b1010010011111010: color_data = 12'b001110100111;
		16'b1010010011111011: color_data = 12'b001110100111;
		16'b1010010011111100: color_data = 12'b001110100111;
		16'b1010010011111101: color_data = 12'b001110100111;
		16'b1010010011111110: color_data = 12'b001110100111;
		16'b1010010011111111: color_data = 12'b001110100111;
		16'b1010010100000000: color_data = 12'b001110100111;
		16'b1010010100000001: color_data = 12'b001110100111;
		16'b1010010100000010: color_data = 12'b001110100111;
		16'b1010010100000011: color_data = 12'b001110100111;
		16'b1010010100000100: color_data = 12'b001110100111;
		16'b1010010100000101: color_data = 12'b001110100111;
		16'b1010010100000110: color_data = 12'b001110100111;
		16'b1010010100000111: color_data = 12'b001110100111;
		16'b1010010100001000: color_data = 12'b001110100111;
		16'b1010010100001001: color_data = 12'b001110100111;
		16'b1010010100001010: color_data = 12'b001110100111;
		16'b1010010100001011: color_data = 12'b001110100111;
		16'b1010010100001100: color_data = 12'b001110100111;
		16'b1010010100001101: color_data = 12'b001110100111;
		16'b1010010100001110: color_data = 12'b001110100111;
		16'b1010010100001111: color_data = 12'b001110100111;
		16'b1010010100010000: color_data = 12'b001110100111;
		16'b1010010100010001: color_data = 12'b001110100111;
		16'b1010010100010010: color_data = 12'b001110100111;
		16'b1010010100010011: color_data = 12'b001110100111;
		16'b1010010100010100: color_data = 12'b001110100111;
		16'b1010010100010101: color_data = 12'b001110100111;
		16'b1010010100010110: color_data = 12'b001110100111;
		16'b1010010100010111: color_data = 12'b001110100111;
		16'b1010010100011000: color_data = 12'b001110100111;
		16'b1010010100011001: color_data = 12'b001110100111;
		16'b1010010100011010: color_data = 12'b001110100111;
		16'b1010010100011011: color_data = 12'b001110100111;
		16'b1010010100011100: color_data = 12'b001110100111;
		16'b1010010100011101: color_data = 12'b001110100111;
		16'b1010010100011110: color_data = 12'b001110100111;
		16'b1010010100011111: color_data = 12'b001110100111;
		16'b1010010100100000: color_data = 12'b001110100111;
		16'b1010010100100001: color_data = 12'b001110100111;
		16'b1010010100100010: color_data = 12'b001110100111;
		16'b1010010100100011: color_data = 12'b001110100111;
		16'b1010010100100100: color_data = 12'b001110100111;
		16'b1010010100100101: color_data = 12'b001110100111;
		16'b1010010100100110: color_data = 12'b001110100111;
		16'b1010010100101101: color_data = 12'b001110100111;
		16'b1010010100101110: color_data = 12'b001110100111;
		16'b1010010100101111: color_data = 12'b001110100111;
		16'b1010010100110000: color_data = 12'b001110100111;
		16'b1010010100110001: color_data = 12'b001110100111;
		16'b1010010100110010: color_data = 12'b001110100111;
		16'b1010010100110011: color_data = 12'b001110100111;
		16'b1010010100110100: color_data = 12'b001110100111;
		16'b1010010100110101: color_data = 12'b001110100111;
		16'b1010010100110110: color_data = 12'b001110100111;
		16'b1010010100110111: color_data = 12'b001110100111;
		16'b1010010100111000: color_data = 12'b001110100111;
		16'b1010010101000101: color_data = 12'b001110100111;
		16'b1010010101000110: color_data = 12'b001110100111;
		16'b1010010101000111: color_data = 12'b001110100111;
		16'b1010010101001000: color_data = 12'b001110100111;
		16'b1010010101001001: color_data = 12'b001110100111;
		16'b1010010101001010: color_data = 12'b001110100111;
		16'b1010010101001011: color_data = 12'b001110100111;
		16'b1010010101001100: color_data = 12'b001110100111;
		16'b1010010101001101: color_data = 12'b001110100111;
		16'b1010010101001110: color_data = 12'b001110100111;
		16'b1010010101001111: color_data = 12'b001110100111;
		16'b1010010101010000: color_data = 12'b001110100111;
		16'b1010010101010001: color_data = 12'b001110100111;
		16'b1010010101011000: color_data = 12'b001110100111;
		16'b1010010101011001: color_data = 12'b001110100111;
		16'b1010010101011010: color_data = 12'b001110100111;
		16'b1010010101011011: color_data = 12'b001110100111;
		16'b1010010101011100: color_data = 12'b001110100111;
		16'b1010010101011101: color_data = 12'b001110100111;
		16'b1010010101011110: color_data = 12'b001110100111;
		16'b1010010101011111: color_data = 12'b001110100111;
		16'b1010010101100000: color_data = 12'b001110100111;
		16'b1010010101100001: color_data = 12'b001110100111;
		16'b1010010101100010: color_data = 12'b001110100111;
		16'b1010010101100011: color_data = 12'b001110100111;
		16'b1010010101100100: color_data = 12'b001110100111;
		16'b1010010101100101: color_data = 12'b001110100111;
		16'b1010010101100110: color_data = 12'b001110100111;
		16'b1010010101100111: color_data = 12'b001110100111;
		16'b1010010101101000: color_data = 12'b001110100111;
		16'b1010010101101001: color_data = 12'b001110100111;
		16'b1010010101101010: color_data = 12'b001110100111;
		16'b1010010101101011: color_data = 12'b001110100111;
		16'b1010010101101100: color_data = 12'b001110100111;
		16'b1010010101101101: color_data = 12'b001110100111;
		16'b1010010101101110: color_data = 12'b001110100111;
		16'b1010010101101111: color_data = 12'b001110100111;
		16'b1010010101110000: color_data = 12'b001110100111;
		16'b1010010101110001: color_data = 12'b001110100111;
		16'b1010010101110010: color_data = 12'b001110100111;
		16'b1010010101110011: color_data = 12'b001110100111;
		16'b1010010101110100: color_data = 12'b001110100111;
		16'b1010010101110101: color_data = 12'b001110100111;
		16'b1010010101110110: color_data = 12'b001110100111;
		16'b1010010101110111: color_data = 12'b001110100111;
		16'b1010010101111000: color_data = 12'b001110100111;
		16'b1010010101111001: color_data = 12'b001110100111;
		16'b1010010101111010: color_data = 12'b001110100111;
		16'b1010010101111011: color_data = 12'b001110100111;
		16'b1010011000000000: color_data = 12'b001110100111;
		16'b1010011000000001: color_data = 12'b001110100111;
		16'b1010011000000010: color_data = 12'b001110100111;
		16'b1010011000000011: color_data = 12'b001110100111;
		16'b1010011000000100: color_data = 12'b001110100111;
		16'b1010011000000101: color_data = 12'b001110100111;
		16'b1010011000000110: color_data = 12'b001110100111;
		16'b1010011000000111: color_data = 12'b001110100111;
		16'b1010011000001000: color_data = 12'b001110100111;
		16'b1010011000001001: color_data = 12'b001110100111;
		16'b1010011000001010: color_data = 12'b001110100111;
		16'b1010011000001011: color_data = 12'b001110100111;
		16'b1010011000001100: color_data = 12'b001110100111;
		16'b1010011000001101: color_data = 12'b001110100111;
		16'b1010011000001110: color_data = 12'b001110100111;
		16'b1010011000001111: color_data = 12'b001110100111;
		16'b1010011000010000: color_data = 12'b001110100111;
		16'b1010011000010001: color_data = 12'b001110100111;
		16'b1010011000010010: color_data = 12'b001110100111;
		16'b1010011000010011: color_data = 12'b001110100111;
		16'b1010011000010100: color_data = 12'b001110100111;
		16'b1010011000010101: color_data = 12'b001110100111;
		16'b1010011000010110: color_data = 12'b001110100111;
		16'b1010011000010111: color_data = 12'b001110100111;
		16'b1010011000011000: color_data = 12'b001110100111;
		16'b1010011000011001: color_data = 12'b001110100111;
		16'b1010011000011010: color_data = 12'b001110100111;
		16'b1010011000011011: color_data = 12'b001110100111;
		16'b1010011000011100: color_data = 12'b001110100111;
		16'b1010011000011101: color_data = 12'b001110100111;
		16'b1010011000011110: color_data = 12'b001110100111;
		16'b1010011000011111: color_data = 12'b001110100111;
		16'b1010011000100000: color_data = 12'b001110100111;
		16'b1010011000100001: color_data = 12'b001110100111;
		16'b1010011000100010: color_data = 12'b001110100111;
		16'b1010011000100011: color_data = 12'b001110100111;
		16'b1010011000100100: color_data = 12'b001110100111;
		16'b1010011000101011: color_data = 12'b001110100111;
		16'b1010011000101100: color_data = 12'b001110100111;
		16'b1010011000101101: color_data = 12'b001110100111;
		16'b1010011000101110: color_data = 12'b001110100111;
		16'b1010011000101111: color_data = 12'b001110100111;
		16'b1010011000110000: color_data = 12'b001110100111;
		16'b1010011000110001: color_data = 12'b001110100111;
		16'b1010011000110010: color_data = 12'b001110100111;
		16'b1010011000110011: color_data = 12'b001110100111;
		16'b1010011000110100: color_data = 12'b001110100111;
		16'b1010011000110101: color_data = 12'b001110100111;
		16'b1010011000110110: color_data = 12'b001110100111;
		16'b1010011000110111: color_data = 12'b001110100111;
		16'b1010011001000100: color_data = 12'b001110100111;
		16'b1010011001000101: color_data = 12'b001110100111;
		16'b1010011001000110: color_data = 12'b001110100111;
		16'b1010011001000111: color_data = 12'b001110100111;
		16'b1010011001001000: color_data = 12'b001110100111;
		16'b1010011001001001: color_data = 12'b001110100111;
		16'b1010011001001010: color_data = 12'b001110100111;
		16'b1010011001001011: color_data = 12'b001110100111;
		16'b1010011001001100: color_data = 12'b001110100111;
		16'b1010011001001101: color_data = 12'b001110100111;
		16'b1010011001001110: color_data = 12'b001110100111;
		16'b1010011001001111: color_data = 12'b001110100111;
		16'b1010011001010110: color_data = 12'b001110100111;
		16'b1010011001010111: color_data = 12'b001110100111;
		16'b1010011001011000: color_data = 12'b001110100111;
		16'b1010011001011001: color_data = 12'b001110100111;
		16'b1010011001011010: color_data = 12'b001110100111;
		16'b1010011001011011: color_data = 12'b001110100111;
		16'b1010011001011100: color_data = 12'b001110100111;
		16'b1010011001011101: color_data = 12'b001110100111;
		16'b1010011001011110: color_data = 12'b001110100111;
		16'b1010011001011111: color_data = 12'b001110100111;
		16'b1010011001100000: color_data = 12'b001110100111;
		16'b1010011001100001: color_data = 12'b001110100111;
		16'b1010011001100010: color_data = 12'b001110100111;
		16'b1010011001100011: color_data = 12'b001110100111;
		16'b1010011001100100: color_data = 12'b001110100111;
		16'b1010011001100101: color_data = 12'b001110100111;
		16'b1010011001100110: color_data = 12'b001110100111;
		16'b1010011001100111: color_data = 12'b001110100111;
		16'b1010011001101000: color_data = 12'b001110100111;
		16'b1010011001101001: color_data = 12'b001110100111;
		16'b1010011001101010: color_data = 12'b001110100111;
		16'b1010011001101011: color_data = 12'b001110100111;
		16'b1010011001101100: color_data = 12'b001110100111;
		16'b1010011001101101: color_data = 12'b001110100111;
		16'b1010011001101110: color_data = 12'b001110100111;
		16'b1010011001110101: color_data = 12'b001110100111;
		16'b1010011001110110: color_data = 12'b001110100111;
		16'b1010011001110111: color_data = 12'b001110100111;
		16'b1010011001111000: color_data = 12'b001110100111;
		16'b1010011001111001: color_data = 12'b001110100111;
		16'b1010011001111010: color_data = 12'b001110100111;
		16'b1010011001111011: color_data = 12'b001110100111;
		16'b1010011001111100: color_data = 12'b001110100111;
		16'b1010011001111101: color_data = 12'b001110100111;
		16'b1010011001111110: color_data = 12'b001110100111;
		16'b1010011001111111: color_data = 12'b001110100111;
		16'b1010011010000000: color_data = 12'b001110100111;
		16'b1010011010001101: color_data = 12'b001110100111;
		16'b1010011010001110: color_data = 12'b001110100111;
		16'b1010011010001111: color_data = 12'b001110100111;
		16'b1010011010010000: color_data = 12'b001110100111;
		16'b1010011010010001: color_data = 12'b001110100111;
		16'b1010011010010010: color_data = 12'b001110100111;
		16'b1010011010010011: color_data = 12'b001110100111;
		16'b1010011010010100: color_data = 12'b001110100111;
		16'b1010011010010101: color_data = 12'b001110100111;
		16'b1010011010010110: color_data = 12'b001110100111;
		16'b1010011010010111: color_data = 12'b001110100111;
		16'b1010011010011000: color_data = 12'b001110100111;
		16'b1010011010011001: color_data = 12'b001110100111;
		16'b1010011010100000: color_data = 12'b001110100111;
		16'b1010011010100001: color_data = 12'b001110100111;
		16'b1010011010100010: color_data = 12'b001110100111;
		16'b1010011010100011: color_data = 12'b001110100111;
		16'b1010011010100100: color_data = 12'b001110100111;
		16'b1010011010100101: color_data = 12'b001110100111;
		16'b1010011010100110: color_data = 12'b001110100111;
		16'b1010011010100111: color_data = 12'b001110100111;
		16'b1010011010101000: color_data = 12'b001110100111;
		16'b1010011010101001: color_data = 12'b001110100111;
		16'b1010011010101010: color_data = 12'b001110100111;
		16'b1010011010101011: color_data = 12'b001110100111;
		16'b1010011010101100: color_data = 12'b001110100111;
		16'b1010011010101101: color_data = 12'b001110100111;
		16'b1010011010101110: color_data = 12'b001110100111;
		16'b1010011010101111: color_data = 12'b001110100111;
		16'b1010011010110000: color_data = 12'b001110100111;
		16'b1010011010110001: color_data = 12'b001110100111;
		16'b1010011010110010: color_data = 12'b001110100111;
		16'b1010011010110011: color_data = 12'b001110100111;
		16'b1010011010110100: color_data = 12'b001110100111;
		16'b1010011010110101: color_data = 12'b001110100111;
		16'b1010011010110110: color_data = 12'b001110100111;
		16'b1010011010110111: color_data = 12'b001110100111;
		16'b1010011010111000: color_data = 12'b001110100111;
		16'b1010011010111001: color_data = 12'b001110100111;
		16'b1010011010111010: color_data = 12'b001110100111;
		16'b1010011010111011: color_data = 12'b001110100111;
		16'b1010011010111100: color_data = 12'b001110100111;
		16'b1010011010111101: color_data = 12'b001110100111;
		16'b1010011010111110: color_data = 12'b001110100111;
		16'b1010011010111111: color_data = 12'b001110100111;
		16'b1010011011000000: color_data = 12'b001110100111;
		16'b1010011011000001: color_data = 12'b001110100111;
		16'b1010011011000010: color_data = 12'b001110100111;
		16'b1010011011000011: color_data = 12'b001110100111;
		16'b1010011011000100: color_data = 12'b001110100111;
		16'b1010011011001011: color_data = 12'b001110100111;
		16'b1010011011001100: color_data = 12'b001110100111;
		16'b1010011011001101: color_data = 12'b001110100111;
		16'b1010011011001110: color_data = 12'b001110100111;
		16'b1010011011001111: color_data = 12'b001110100111;
		16'b1010011011010000: color_data = 12'b001110100111;
		16'b1010011011010001: color_data = 12'b001110100111;
		16'b1010011011010010: color_data = 12'b001110100111;
		16'b1010011011010011: color_data = 12'b001110100111;
		16'b1010011011010100: color_data = 12'b001110100111;
		16'b1010011011010101: color_data = 12'b001110100111;
		16'b1010011011010110: color_data = 12'b001110100111;
		16'b1010011011110110: color_data = 12'b001110100111;
		16'b1010011011110111: color_data = 12'b001110100111;
		16'b1010011011111000: color_data = 12'b001110100111;
		16'b1010011011111001: color_data = 12'b001110100111;
		16'b1010011011111010: color_data = 12'b001110100111;
		16'b1010011011111011: color_data = 12'b001110100111;
		16'b1010011011111100: color_data = 12'b001110100111;
		16'b1010011011111101: color_data = 12'b001110100111;
		16'b1010011011111110: color_data = 12'b001110100111;
		16'b1010011011111111: color_data = 12'b001110100111;
		16'b1010011100000000: color_data = 12'b001110100111;
		16'b1010011100000001: color_data = 12'b001110100111;
		16'b1010011100000010: color_data = 12'b001110100111;
		16'b1010011100000011: color_data = 12'b001110100111;
		16'b1010011100000100: color_data = 12'b001110100111;
		16'b1010011100000101: color_data = 12'b001110100111;
		16'b1010011100000110: color_data = 12'b001110100111;
		16'b1010011100000111: color_data = 12'b001110100111;
		16'b1010011100001000: color_data = 12'b001110100111;
		16'b1010011100001001: color_data = 12'b001110100111;
		16'b1010011100001010: color_data = 12'b001110100111;
		16'b1010011100001011: color_data = 12'b001110100111;
		16'b1010011100001100: color_data = 12'b001110100111;
		16'b1010011100001101: color_data = 12'b001110100111;
		16'b1010011100001110: color_data = 12'b001110100111;
		16'b1010011100001111: color_data = 12'b001110100111;
		16'b1010011100010000: color_data = 12'b001110100111;
		16'b1010011100010001: color_data = 12'b001110100111;
		16'b1010011100010010: color_data = 12'b001110100111;
		16'b1010011100010011: color_data = 12'b001110100111;
		16'b1010011100010100: color_data = 12'b001110100111;
		16'b1010011100010101: color_data = 12'b001110100111;
		16'b1010011100010110: color_data = 12'b001110100111;
		16'b1010011100010111: color_data = 12'b001110100111;
		16'b1010011100011000: color_data = 12'b001110100111;
		16'b1010011100011001: color_data = 12'b001110100111;
		16'b1010011100011010: color_data = 12'b001110100111;
		16'b1010011100011011: color_data = 12'b001110100111;
		16'b1010011100011100: color_data = 12'b001110100111;
		16'b1010011100011101: color_data = 12'b001110100111;
		16'b1010011100011110: color_data = 12'b001110100111;
		16'b1010011100011111: color_data = 12'b001110100111;
		16'b1010011100100000: color_data = 12'b001110100111;
		16'b1010011100100001: color_data = 12'b001110100111;
		16'b1010011100100010: color_data = 12'b001110100111;
		16'b1010011100100011: color_data = 12'b001110100111;
		16'b1010011100100100: color_data = 12'b001110100111;
		16'b1010011100100101: color_data = 12'b001110100111;
		16'b1010011100100110: color_data = 12'b001110100111;
		16'b1010011100101101: color_data = 12'b001110100111;
		16'b1010011100101110: color_data = 12'b001110100111;
		16'b1010011100101111: color_data = 12'b001110100111;
		16'b1010011100110000: color_data = 12'b001110100111;
		16'b1010011100110001: color_data = 12'b001110100111;
		16'b1010011100110010: color_data = 12'b001110100111;
		16'b1010011100110011: color_data = 12'b001110100111;
		16'b1010011100110100: color_data = 12'b001110100111;
		16'b1010011100110101: color_data = 12'b001110100111;
		16'b1010011100110110: color_data = 12'b001110100111;
		16'b1010011100110111: color_data = 12'b001110100111;
		16'b1010011100111000: color_data = 12'b001110100111;
		16'b1010011101000101: color_data = 12'b001110100111;
		16'b1010011101000110: color_data = 12'b001110100111;
		16'b1010011101000111: color_data = 12'b001110100111;
		16'b1010011101001000: color_data = 12'b001110100111;
		16'b1010011101001001: color_data = 12'b001110100111;
		16'b1010011101001010: color_data = 12'b001110100111;
		16'b1010011101001011: color_data = 12'b001110100111;
		16'b1010011101001100: color_data = 12'b001110100111;
		16'b1010011101001101: color_data = 12'b001110100111;
		16'b1010011101001110: color_data = 12'b001110100111;
		16'b1010011101001111: color_data = 12'b001110100111;
		16'b1010011101010000: color_data = 12'b001110100111;
		16'b1010011101010001: color_data = 12'b001110100111;
		16'b1010011101011000: color_data = 12'b001110100111;
		16'b1010011101011001: color_data = 12'b001110100111;
		16'b1010011101011010: color_data = 12'b001110100111;
		16'b1010011101011011: color_data = 12'b001110100111;
		16'b1010011101011100: color_data = 12'b001110100111;
		16'b1010011101011101: color_data = 12'b001110100111;
		16'b1010011101011110: color_data = 12'b001110100111;
		16'b1010011101011111: color_data = 12'b001110100111;
		16'b1010011101100000: color_data = 12'b001110100111;
		16'b1010011101100001: color_data = 12'b001110100111;
		16'b1010011101100010: color_data = 12'b001110100111;
		16'b1010011101100011: color_data = 12'b001110100111;
		16'b1010011101100100: color_data = 12'b001110100111;
		16'b1010011101100101: color_data = 12'b001110100111;
		16'b1010011101100110: color_data = 12'b001110100111;
		16'b1010011101100111: color_data = 12'b001110100111;
		16'b1010011101101000: color_data = 12'b001110100111;
		16'b1010011101101001: color_data = 12'b001110100111;
		16'b1010011101101010: color_data = 12'b001110100111;
		16'b1010011101101011: color_data = 12'b001110100111;
		16'b1010011101101100: color_data = 12'b001110100111;
		16'b1010011101101101: color_data = 12'b001110100111;
		16'b1010011101101110: color_data = 12'b001110100111;
		16'b1010011101101111: color_data = 12'b001110100111;
		16'b1010011101110000: color_data = 12'b001110100111;
		16'b1010011101110001: color_data = 12'b001110100111;
		16'b1010011101110010: color_data = 12'b001110100111;
		16'b1010011101110011: color_data = 12'b001110100111;
		16'b1010011101110100: color_data = 12'b001110100111;
		16'b1010011101110101: color_data = 12'b001110100111;
		16'b1010011101110110: color_data = 12'b001110100111;
		16'b1010011101110111: color_data = 12'b001110100111;
		16'b1010011101111000: color_data = 12'b001110100111;
		16'b1010011101111001: color_data = 12'b001110100111;
		16'b1010011101111010: color_data = 12'b001110100111;
		16'b1010011101111011: color_data = 12'b001110100111;
		16'b1010100000000000: color_data = 12'b001110100111;
		16'b1010100000000001: color_data = 12'b001110100111;
		16'b1010100000000010: color_data = 12'b001110100111;
		16'b1010100000000011: color_data = 12'b001110100111;
		16'b1010100000000100: color_data = 12'b001110100111;
		16'b1010100000000101: color_data = 12'b001110100111;
		16'b1010100000000110: color_data = 12'b001110100111;
		16'b1010100000000111: color_data = 12'b001110100111;
		16'b1010100000001000: color_data = 12'b001110100111;
		16'b1010100000001001: color_data = 12'b001110100111;
		16'b1010100000001010: color_data = 12'b001110100111;
		16'b1010100000001011: color_data = 12'b001110100111;
		16'b1010100000001100: color_data = 12'b001110100111;
		16'b1010100000001101: color_data = 12'b001110100111;
		16'b1010100000001110: color_data = 12'b001110100111;
		16'b1010100000001111: color_data = 12'b001110100111;
		16'b1010100000010000: color_data = 12'b001110100111;
		16'b1010100000010001: color_data = 12'b001110100111;
		16'b1010100000010010: color_data = 12'b001110100111;
		16'b1010100000010011: color_data = 12'b001110100111;
		16'b1010100000010100: color_data = 12'b001110100111;
		16'b1010100000010101: color_data = 12'b001110100111;
		16'b1010100000010110: color_data = 12'b001110100111;
		16'b1010100000010111: color_data = 12'b001110100111;
		16'b1010100000011000: color_data = 12'b001110100111;
		16'b1010100000011001: color_data = 12'b001110100111;
		16'b1010100000011010: color_data = 12'b001110100111;
		16'b1010100000011011: color_data = 12'b001110100111;
		16'b1010100000011100: color_data = 12'b001110100111;
		16'b1010100000011101: color_data = 12'b001110100111;
		16'b1010100000011110: color_data = 12'b001110100111;
		16'b1010100000011111: color_data = 12'b001110100111;
		16'b1010100000100000: color_data = 12'b001110100111;
		16'b1010100000100001: color_data = 12'b001110100111;
		16'b1010100000100010: color_data = 12'b001110100111;
		16'b1010100000100011: color_data = 12'b001110100111;
		16'b1010100000100100: color_data = 12'b001110100111;
		16'b1010100000101011: color_data = 12'b001110100111;
		16'b1010100000101100: color_data = 12'b001110100111;
		16'b1010100000101101: color_data = 12'b001110100111;
		16'b1010100000101110: color_data = 12'b001110100111;
		16'b1010100000101111: color_data = 12'b001110100111;
		16'b1010100000110000: color_data = 12'b001110100111;
		16'b1010100000110001: color_data = 12'b001110100111;
		16'b1010100000110010: color_data = 12'b001110100111;
		16'b1010100000110011: color_data = 12'b001110100111;
		16'b1010100000110100: color_data = 12'b001110100111;
		16'b1010100000110101: color_data = 12'b001110100111;
		16'b1010100000110110: color_data = 12'b001110100111;
		16'b1010100000110111: color_data = 12'b001110100111;
		16'b1010100001000100: color_data = 12'b001110100111;
		16'b1010100001000101: color_data = 12'b001110100111;
		16'b1010100001000110: color_data = 12'b001110100111;
		16'b1010100001000111: color_data = 12'b001110100111;
		16'b1010100001001000: color_data = 12'b001110100111;
		16'b1010100001001001: color_data = 12'b001110100111;
		16'b1010100001001010: color_data = 12'b001110100111;
		16'b1010100001001011: color_data = 12'b001110100111;
		16'b1010100001001100: color_data = 12'b001110100111;
		16'b1010100001001101: color_data = 12'b001110100111;
		16'b1010100001001110: color_data = 12'b001110100111;
		16'b1010100001001111: color_data = 12'b001110100111;
		16'b1010100001010110: color_data = 12'b001110100111;
		16'b1010100001010111: color_data = 12'b001110100111;
		16'b1010100001011000: color_data = 12'b001110100111;
		16'b1010100001011001: color_data = 12'b001110100111;
		16'b1010100001011010: color_data = 12'b001110100111;
		16'b1010100001011011: color_data = 12'b001110100111;
		16'b1010100001011100: color_data = 12'b001110100111;
		16'b1010100001011101: color_data = 12'b001110100111;
		16'b1010100001011110: color_data = 12'b001110100111;
		16'b1010100001011111: color_data = 12'b001110100111;
		16'b1010100001100000: color_data = 12'b001110100111;
		16'b1010100001100001: color_data = 12'b001110100111;
		16'b1010100001100010: color_data = 12'b001110100111;
		16'b1010100001100011: color_data = 12'b001110100111;
		16'b1010100001100100: color_data = 12'b001110100111;
		16'b1010100001100101: color_data = 12'b001110100111;
		16'b1010100001100110: color_data = 12'b001110100111;
		16'b1010100001100111: color_data = 12'b001110100111;
		16'b1010100001101000: color_data = 12'b001110100111;
		16'b1010100001101001: color_data = 12'b001110100111;
		16'b1010100001101010: color_data = 12'b001110100111;
		16'b1010100001101011: color_data = 12'b001110100111;
		16'b1010100001101100: color_data = 12'b001110100111;
		16'b1010100001101101: color_data = 12'b001110100111;
		16'b1010100001101110: color_data = 12'b001110100111;
		16'b1010100001110101: color_data = 12'b001110100111;
		16'b1010100001110110: color_data = 12'b001110100111;
		16'b1010100001110111: color_data = 12'b001110100111;
		16'b1010100001111000: color_data = 12'b001110100111;
		16'b1010100001111001: color_data = 12'b001110100111;
		16'b1010100001111010: color_data = 12'b001110100111;
		16'b1010100001111011: color_data = 12'b001110100111;
		16'b1010100001111100: color_data = 12'b001110100111;
		16'b1010100001111101: color_data = 12'b001110100111;
		16'b1010100001111110: color_data = 12'b001110100111;
		16'b1010100001111111: color_data = 12'b001110100111;
		16'b1010100010000000: color_data = 12'b001110100111;
		16'b1010100010001101: color_data = 12'b001110100111;
		16'b1010100010001110: color_data = 12'b001110100111;
		16'b1010100010001111: color_data = 12'b001110100111;
		16'b1010100010010000: color_data = 12'b001110100111;
		16'b1010100010010001: color_data = 12'b001110100111;
		16'b1010100010010010: color_data = 12'b001110100111;
		16'b1010100010010011: color_data = 12'b001110100111;
		16'b1010100010010100: color_data = 12'b001110100111;
		16'b1010100010010101: color_data = 12'b001110100111;
		16'b1010100010010110: color_data = 12'b001110100111;
		16'b1010100010010111: color_data = 12'b001110100111;
		16'b1010100010011000: color_data = 12'b001110100111;
		16'b1010100010011001: color_data = 12'b001110100111;
		16'b1010100010100000: color_data = 12'b001110100111;
		16'b1010100010100001: color_data = 12'b001110100111;
		16'b1010100010100010: color_data = 12'b001110100111;
		16'b1010100010100011: color_data = 12'b001110100111;
		16'b1010100010100100: color_data = 12'b001110100111;
		16'b1010100010100101: color_data = 12'b001110100111;
		16'b1010100010100110: color_data = 12'b001110100111;
		16'b1010100010100111: color_data = 12'b001110100111;
		16'b1010100010101000: color_data = 12'b001110100111;
		16'b1010100010101001: color_data = 12'b001110100111;
		16'b1010100010101010: color_data = 12'b001110100111;
		16'b1010100010101011: color_data = 12'b001110100111;
		16'b1010100010101100: color_data = 12'b001110100111;
		16'b1010100010101101: color_data = 12'b001110100111;
		16'b1010100010101110: color_data = 12'b001110100111;
		16'b1010100010101111: color_data = 12'b001110100111;
		16'b1010100010110000: color_data = 12'b001110100111;
		16'b1010100010110001: color_data = 12'b001110100111;
		16'b1010100010110010: color_data = 12'b001110100111;
		16'b1010100010110011: color_data = 12'b001110100111;
		16'b1010100010110100: color_data = 12'b001110100111;
		16'b1010100010110101: color_data = 12'b001110100111;
		16'b1010100010110110: color_data = 12'b001110100111;
		16'b1010100010110111: color_data = 12'b001110100111;
		16'b1010100010111000: color_data = 12'b001110100111;
		16'b1010100010111001: color_data = 12'b001110100111;
		16'b1010100010111010: color_data = 12'b001110100111;
		16'b1010100010111011: color_data = 12'b001110100111;
		16'b1010100010111100: color_data = 12'b001110100111;
		16'b1010100010111101: color_data = 12'b001110100111;
		16'b1010100010111110: color_data = 12'b001110100111;
		16'b1010100010111111: color_data = 12'b001110100111;
		16'b1010100011000000: color_data = 12'b001110100111;
		16'b1010100011000001: color_data = 12'b001110100111;
		16'b1010100011000010: color_data = 12'b001110100111;
		16'b1010100011000011: color_data = 12'b001110100111;
		16'b1010100011000100: color_data = 12'b001110100111;
		16'b1010100011001011: color_data = 12'b001110100111;
		16'b1010100011001100: color_data = 12'b001110100111;
		16'b1010100011001101: color_data = 12'b001110100111;
		16'b1010100011001110: color_data = 12'b001110100111;
		16'b1010100011001111: color_data = 12'b001110100111;
		16'b1010100011010000: color_data = 12'b001110100111;
		16'b1010100011010001: color_data = 12'b001110100111;
		16'b1010100011010010: color_data = 12'b001110100111;
		16'b1010100011010011: color_data = 12'b001110100111;
		16'b1010100011010100: color_data = 12'b001110100111;
		16'b1010100011010101: color_data = 12'b001110100111;
		16'b1010100011010110: color_data = 12'b001110100111;
		16'b1010100011110110: color_data = 12'b001110100111;
		16'b1010100011110111: color_data = 12'b001110100111;
		16'b1010100011111000: color_data = 12'b001110100111;
		16'b1010100011111001: color_data = 12'b001110100111;
		16'b1010100011111010: color_data = 12'b001110100111;
		16'b1010100011111011: color_data = 12'b001110100111;
		16'b1010100011111100: color_data = 12'b001110100111;
		16'b1010100011111101: color_data = 12'b001110100111;
		16'b1010100011111110: color_data = 12'b001110100111;
		16'b1010100011111111: color_data = 12'b001110100111;
		16'b1010100100000000: color_data = 12'b001110100111;
		16'b1010100100000001: color_data = 12'b001110100111;
		16'b1010100100000010: color_data = 12'b001110100111;
		16'b1010100100000011: color_data = 12'b001110100111;
		16'b1010100100000100: color_data = 12'b001110100111;
		16'b1010100100000101: color_data = 12'b001110100111;
		16'b1010100100000110: color_data = 12'b001110100111;
		16'b1010100100000111: color_data = 12'b001110100111;
		16'b1010100100001000: color_data = 12'b001110100111;
		16'b1010100100001001: color_data = 12'b001110100111;
		16'b1010100100001010: color_data = 12'b001110100111;
		16'b1010100100001011: color_data = 12'b001110100111;
		16'b1010100100001100: color_data = 12'b001110100111;
		16'b1010100100001101: color_data = 12'b001110100111;
		16'b1010100100001110: color_data = 12'b001110100111;
		16'b1010100100001111: color_data = 12'b001110100111;
		16'b1010100100010000: color_data = 12'b001110100111;
		16'b1010100100010001: color_data = 12'b001110100111;
		16'b1010100100010010: color_data = 12'b001110100111;
		16'b1010100100010011: color_data = 12'b001110100111;
		16'b1010100100010100: color_data = 12'b001110100111;
		16'b1010100100010101: color_data = 12'b001110100111;
		16'b1010100100010110: color_data = 12'b001110100111;
		16'b1010100100010111: color_data = 12'b001110100111;
		16'b1010100100011000: color_data = 12'b001110100111;
		16'b1010100100011001: color_data = 12'b001110100111;
		16'b1010100100011010: color_data = 12'b001110100111;
		16'b1010100100011011: color_data = 12'b001110100111;
		16'b1010100100011100: color_data = 12'b001110100111;
		16'b1010100100011101: color_data = 12'b001110100111;
		16'b1010100100011110: color_data = 12'b001110100111;
		16'b1010100100011111: color_data = 12'b001110100111;
		16'b1010100100100000: color_data = 12'b001110100111;
		16'b1010100100100001: color_data = 12'b001110100111;
		16'b1010100100100010: color_data = 12'b001110100111;
		16'b1010100100100011: color_data = 12'b001110100111;
		16'b1010100100100100: color_data = 12'b001110100111;
		16'b1010100100100101: color_data = 12'b001110100111;
		16'b1010100100100110: color_data = 12'b001110100111;
		16'b1010100100101101: color_data = 12'b001110100111;
		16'b1010100100101110: color_data = 12'b001110100111;
		16'b1010100100101111: color_data = 12'b001110100111;
		16'b1010100100110000: color_data = 12'b001110100111;
		16'b1010100100110001: color_data = 12'b001110100111;
		16'b1010100100110010: color_data = 12'b001110100111;
		16'b1010100100110011: color_data = 12'b001110100111;
		16'b1010100100110100: color_data = 12'b001110100111;
		16'b1010100100110101: color_data = 12'b001110100111;
		16'b1010100100110110: color_data = 12'b001110100111;
		16'b1010100100110111: color_data = 12'b001110100111;
		16'b1010100100111000: color_data = 12'b001110100111;
		16'b1010100101000101: color_data = 12'b001110100111;
		16'b1010100101000110: color_data = 12'b001110100111;
		16'b1010100101000111: color_data = 12'b001110100111;
		16'b1010100101001000: color_data = 12'b001110100111;
		16'b1010100101001001: color_data = 12'b001110100111;
		16'b1010100101001010: color_data = 12'b001110100111;
		16'b1010100101001011: color_data = 12'b001110100111;
		16'b1010100101001100: color_data = 12'b001110100111;
		16'b1010100101001101: color_data = 12'b001110100111;
		16'b1010100101001110: color_data = 12'b001110100111;
		16'b1010100101001111: color_data = 12'b001110100111;
		16'b1010100101010000: color_data = 12'b001110100111;
		16'b1010100101010001: color_data = 12'b001110100111;
		16'b1010100101011000: color_data = 12'b001110100111;
		16'b1010100101011001: color_data = 12'b001110100111;
		16'b1010100101011010: color_data = 12'b001110100111;
		16'b1010100101011011: color_data = 12'b001110100111;
		16'b1010100101011100: color_data = 12'b001110100111;
		16'b1010100101011101: color_data = 12'b001110100111;
		16'b1010100101011110: color_data = 12'b001110100111;
		16'b1010100101011111: color_data = 12'b001110100111;
		16'b1010100101100000: color_data = 12'b001110100111;
		16'b1010100101100001: color_data = 12'b001110100111;
		16'b1010100101100010: color_data = 12'b001110100111;
		16'b1010100101100011: color_data = 12'b001110100111;
		16'b1010100101100100: color_data = 12'b001110100111;
		16'b1010100101100101: color_data = 12'b001110100111;
		16'b1010100101100110: color_data = 12'b001110100111;
		16'b1010100101100111: color_data = 12'b001110100111;
		16'b1010100101101000: color_data = 12'b001110100111;
		16'b1010100101101001: color_data = 12'b001110100111;
		16'b1010100101101010: color_data = 12'b001110100111;
		16'b1010100101101011: color_data = 12'b001110100111;
		16'b1010100101101100: color_data = 12'b001110100111;
		16'b1010100101101101: color_data = 12'b001110100111;
		16'b1010100101101110: color_data = 12'b001110100111;
		16'b1010100101101111: color_data = 12'b001110100111;
		16'b1010100101110000: color_data = 12'b001110100111;
		16'b1010100101110001: color_data = 12'b001110100111;
		16'b1010100101110010: color_data = 12'b001110100111;
		16'b1010100101110011: color_data = 12'b001110100111;
		16'b1010100101110100: color_data = 12'b001110100111;
		16'b1010100101110101: color_data = 12'b001110100111;
		16'b1010100101110110: color_data = 12'b001110100111;
		16'b1010100101110111: color_data = 12'b001110100111;
		16'b1010100101111000: color_data = 12'b001110100111;
		16'b1010100101111001: color_data = 12'b001110100111;
		16'b1010100101111010: color_data = 12'b001110100111;
		16'b1010100101111011: color_data = 12'b001110100111;
		16'b1010101000000000: color_data = 12'b001110100111;
		16'b1010101000000001: color_data = 12'b001110100111;
		16'b1010101000000010: color_data = 12'b001110100111;
		16'b1010101000000011: color_data = 12'b001110100111;
		16'b1010101000000100: color_data = 12'b001110100111;
		16'b1010101000000101: color_data = 12'b001110100111;
		16'b1010101000000110: color_data = 12'b001110100111;
		16'b1010101000000111: color_data = 12'b001110100111;
		16'b1010101000001000: color_data = 12'b001110100111;
		16'b1010101000001001: color_data = 12'b001110100111;
		16'b1010101000001010: color_data = 12'b001110100111;
		16'b1010101000001011: color_data = 12'b001110100111;
		16'b1010101000001100: color_data = 12'b001110100111;
		16'b1010101000001101: color_data = 12'b001110100111;
		16'b1010101000001110: color_data = 12'b001110100111;
		16'b1010101000001111: color_data = 12'b001110100111;
		16'b1010101000010000: color_data = 12'b001110100111;
		16'b1010101000010001: color_data = 12'b001110100111;
		16'b1010101000010010: color_data = 12'b001110100111;
		16'b1010101000010011: color_data = 12'b001110100111;
		16'b1010101000010100: color_data = 12'b001110100111;
		16'b1010101000010101: color_data = 12'b001110100111;
		16'b1010101000010110: color_data = 12'b001110100111;
		16'b1010101000010111: color_data = 12'b001110100111;
		16'b1010101000011000: color_data = 12'b001110100111;
		16'b1010101000011001: color_data = 12'b001110100111;
		16'b1010101000011010: color_data = 12'b001110100111;
		16'b1010101000011011: color_data = 12'b001110100111;
		16'b1010101000011100: color_data = 12'b001110100111;
		16'b1010101000011101: color_data = 12'b001110100111;
		16'b1010101000011110: color_data = 12'b001110100111;
		16'b1010101000011111: color_data = 12'b001110100111;
		16'b1010101000100000: color_data = 12'b001110100111;
		16'b1010101000100001: color_data = 12'b001110100111;
		16'b1010101000100010: color_data = 12'b001110100111;
		16'b1010101000100011: color_data = 12'b001110100111;
		16'b1010101000100100: color_data = 12'b001110100111;
		16'b1010101000101011: color_data = 12'b001110100111;
		16'b1010101000101100: color_data = 12'b001110100111;
		16'b1010101000101101: color_data = 12'b001110100111;
		16'b1010101000101110: color_data = 12'b001110100111;
		16'b1010101000101111: color_data = 12'b001110100111;
		16'b1010101000110000: color_data = 12'b001110100111;
		16'b1010101000110001: color_data = 12'b001110100111;
		16'b1010101000110010: color_data = 12'b001110100111;
		16'b1010101000110011: color_data = 12'b001110100111;
		16'b1010101000110100: color_data = 12'b001110100111;
		16'b1010101000110101: color_data = 12'b001110100111;
		16'b1010101000110110: color_data = 12'b001110100111;
		16'b1010101000110111: color_data = 12'b001110100111;
		16'b1010101001000100: color_data = 12'b001110100111;
		16'b1010101001000101: color_data = 12'b001110100111;
		16'b1010101001000110: color_data = 12'b001110100111;
		16'b1010101001000111: color_data = 12'b001110100111;
		16'b1010101001001000: color_data = 12'b001110100111;
		16'b1010101001001001: color_data = 12'b001110100111;
		16'b1010101001001010: color_data = 12'b001110100111;
		16'b1010101001001011: color_data = 12'b001110100111;
		16'b1010101001001100: color_data = 12'b001110100111;
		16'b1010101001001101: color_data = 12'b001110100111;
		16'b1010101001001110: color_data = 12'b001110100111;
		16'b1010101001001111: color_data = 12'b001110100111;
		16'b1010101001010110: color_data = 12'b001110100111;
		16'b1010101001010111: color_data = 12'b001110100111;
		16'b1010101001011000: color_data = 12'b001110100111;
		16'b1010101001011001: color_data = 12'b001110100111;
		16'b1010101001011010: color_data = 12'b001110100111;
		16'b1010101001011011: color_data = 12'b001110100111;
		16'b1010101001011100: color_data = 12'b001110100111;
		16'b1010101001011101: color_data = 12'b001110100111;
		16'b1010101001011110: color_data = 12'b001110100111;
		16'b1010101001011111: color_data = 12'b001110100111;
		16'b1010101001100000: color_data = 12'b001110100111;
		16'b1010101001100001: color_data = 12'b001110100111;
		16'b1010101001100010: color_data = 12'b001110100111;
		16'b1010101001100011: color_data = 12'b001110100111;
		16'b1010101001100100: color_data = 12'b001110100111;
		16'b1010101001100101: color_data = 12'b001110100111;
		16'b1010101001100110: color_data = 12'b001110100111;
		16'b1010101001100111: color_data = 12'b001110100111;
		16'b1010101001101000: color_data = 12'b001110100111;
		16'b1010101001101001: color_data = 12'b001110100111;
		16'b1010101001101010: color_data = 12'b001110100111;
		16'b1010101001101011: color_data = 12'b001110100111;
		16'b1010101001101100: color_data = 12'b001110100111;
		16'b1010101001101101: color_data = 12'b001110100111;
		16'b1010101001101110: color_data = 12'b001110100111;
		16'b1010101001110101: color_data = 12'b001110100111;
		16'b1010101001110110: color_data = 12'b001110100111;
		16'b1010101001110111: color_data = 12'b001110100111;
		16'b1010101001111000: color_data = 12'b001110100111;
		16'b1010101001111001: color_data = 12'b001110100111;
		16'b1010101001111010: color_data = 12'b001110100111;
		16'b1010101001111011: color_data = 12'b001110100111;
		16'b1010101001111100: color_data = 12'b001110100111;
		16'b1010101001111101: color_data = 12'b001110100111;
		16'b1010101001111110: color_data = 12'b001110100111;
		16'b1010101001111111: color_data = 12'b001110100111;
		16'b1010101010000000: color_data = 12'b001110100111;
		16'b1010101010001101: color_data = 12'b001110100111;
		16'b1010101010001110: color_data = 12'b001110100111;
		16'b1010101010001111: color_data = 12'b001110100111;
		16'b1010101010010000: color_data = 12'b001110100111;
		16'b1010101010010001: color_data = 12'b001110100111;
		16'b1010101010010010: color_data = 12'b001110100111;
		16'b1010101010010011: color_data = 12'b001110100111;
		16'b1010101010010100: color_data = 12'b001110100111;
		16'b1010101010010101: color_data = 12'b001110100111;
		16'b1010101010010110: color_data = 12'b001110100111;
		16'b1010101010010111: color_data = 12'b001110100111;
		16'b1010101010011000: color_data = 12'b001110100111;
		16'b1010101010011001: color_data = 12'b001110100111;
		16'b1010101010100000: color_data = 12'b001110100111;
		16'b1010101010100001: color_data = 12'b001110100111;
		16'b1010101010100010: color_data = 12'b001110100111;
		16'b1010101010100011: color_data = 12'b001110100111;
		16'b1010101010100100: color_data = 12'b001110100111;
		16'b1010101010100101: color_data = 12'b001110100111;
		16'b1010101010100110: color_data = 12'b001110100111;
		16'b1010101010100111: color_data = 12'b001110100111;
		16'b1010101010101000: color_data = 12'b001110100111;
		16'b1010101010101001: color_data = 12'b001110100111;
		16'b1010101010101010: color_data = 12'b001110100111;
		16'b1010101010101011: color_data = 12'b001110100111;
		16'b1010101010101100: color_data = 12'b001110100111;
		16'b1010101010101101: color_data = 12'b001110100111;
		16'b1010101010101110: color_data = 12'b001110100111;
		16'b1010101010101111: color_data = 12'b001110100111;
		16'b1010101010110000: color_data = 12'b001110100111;
		16'b1010101010110001: color_data = 12'b001110100111;
		16'b1010101010110010: color_data = 12'b001110100111;
		16'b1010101010110011: color_data = 12'b001110100111;
		16'b1010101010110100: color_data = 12'b001110100111;
		16'b1010101010110101: color_data = 12'b001110100111;
		16'b1010101010110110: color_data = 12'b001110100111;
		16'b1010101010110111: color_data = 12'b001110100111;
		16'b1010101010111000: color_data = 12'b001110100111;
		16'b1010101010111001: color_data = 12'b001110100111;
		16'b1010101010111010: color_data = 12'b001110100111;
		16'b1010101010111011: color_data = 12'b001110100111;
		16'b1010101010111100: color_data = 12'b001110100111;
		16'b1010101010111101: color_data = 12'b001110100111;
		16'b1010101010111110: color_data = 12'b001110100111;
		16'b1010101010111111: color_data = 12'b001110100111;
		16'b1010101011000000: color_data = 12'b001110100111;
		16'b1010101011000001: color_data = 12'b001110100111;
		16'b1010101011000010: color_data = 12'b001110100111;
		16'b1010101011000011: color_data = 12'b001110100111;
		16'b1010101011000100: color_data = 12'b001110100111;
		16'b1010101011001011: color_data = 12'b001110100111;
		16'b1010101011001100: color_data = 12'b001110100111;
		16'b1010101011001101: color_data = 12'b001110100111;
		16'b1010101011001110: color_data = 12'b001110100111;
		16'b1010101011001111: color_data = 12'b001110100111;
		16'b1010101011010000: color_data = 12'b001110100111;
		16'b1010101011010001: color_data = 12'b001110100111;
		16'b1010101011010010: color_data = 12'b001110100111;
		16'b1010101011010011: color_data = 12'b001110100111;
		16'b1010101011010100: color_data = 12'b001110100111;
		16'b1010101011010101: color_data = 12'b001110100111;
		16'b1010101011010110: color_data = 12'b001110100111;
		16'b1010101011110110: color_data = 12'b001110100111;
		16'b1010101011110111: color_data = 12'b001110100111;
		16'b1010101011111000: color_data = 12'b001110100111;
		16'b1010101011111001: color_data = 12'b001110100111;
		16'b1010101011111010: color_data = 12'b001110100111;
		16'b1010101011111011: color_data = 12'b001110100111;
		16'b1010101011111100: color_data = 12'b001110100111;
		16'b1010101011111101: color_data = 12'b001110100111;
		16'b1010101011111110: color_data = 12'b001110100111;
		16'b1010101011111111: color_data = 12'b001110100111;
		16'b1010101100000000: color_data = 12'b001110100111;
		16'b1010101100000001: color_data = 12'b001110100111;
		16'b1010101100000010: color_data = 12'b001110100111;
		16'b1010101100000011: color_data = 12'b001110100111;
		16'b1010101100000100: color_data = 12'b001110100111;
		16'b1010101100000101: color_data = 12'b001110100111;
		16'b1010101100000110: color_data = 12'b001110100111;
		16'b1010101100000111: color_data = 12'b001110100111;
		16'b1010101100001000: color_data = 12'b001110100111;
		16'b1010101100001001: color_data = 12'b001110100111;
		16'b1010101100001010: color_data = 12'b001110100111;
		16'b1010101100001011: color_data = 12'b001110100111;
		16'b1010101100001100: color_data = 12'b001110100111;
		16'b1010101100001101: color_data = 12'b001110100111;
		16'b1010101100001110: color_data = 12'b001110100111;
		16'b1010101100001111: color_data = 12'b001110100111;
		16'b1010101100010000: color_data = 12'b001110100111;
		16'b1010101100010001: color_data = 12'b001110100111;
		16'b1010101100010010: color_data = 12'b001110100111;
		16'b1010101100010011: color_data = 12'b001110100111;
		16'b1010101100010100: color_data = 12'b001110100111;
		16'b1010101100010101: color_data = 12'b001110100111;
		16'b1010101100010110: color_data = 12'b001110100111;
		16'b1010101100010111: color_data = 12'b001110100111;
		16'b1010101100011000: color_data = 12'b001110100111;
		16'b1010101100011001: color_data = 12'b001110100111;
		16'b1010101100011010: color_data = 12'b001110100111;
		16'b1010101100011011: color_data = 12'b001110100111;
		16'b1010101100011100: color_data = 12'b001110100111;
		16'b1010101100011101: color_data = 12'b001110100111;
		16'b1010101100011110: color_data = 12'b001110100111;
		16'b1010101100011111: color_data = 12'b001110100111;
		16'b1010101100100000: color_data = 12'b001110100111;
		16'b1010101100100001: color_data = 12'b001110100111;
		16'b1010101100100010: color_data = 12'b001110100111;
		16'b1010101100100011: color_data = 12'b001110100111;
		16'b1010101100100100: color_data = 12'b001110100111;
		16'b1010101100100101: color_data = 12'b001110100111;
		16'b1010101100100110: color_data = 12'b001110100111;
		16'b1010101100101101: color_data = 12'b001110100111;
		16'b1010101100101110: color_data = 12'b001110100111;
		16'b1010101100101111: color_data = 12'b001110100111;
		16'b1010101100110000: color_data = 12'b001110100111;
		16'b1010101100110001: color_data = 12'b001110100111;
		16'b1010101100110010: color_data = 12'b001110100111;
		16'b1010101100110011: color_data = 12'b001110100111;
		16'b1010101100110100: color_data = 12'b001110100111;
		16'b1010101100110101: color_data = 12'b001110100111;
		16'b1010101100110110: color_data = 12'b001110100111;
		16'b1010101100110111: color_data = 12'b001110100111;
		16'b1010101100111000: color_data = 12'b001110100111;
		16'b1010101101000101: color_data = 12'b001110100111;
		16'b1010101101000110: color_data = 12'b001110100111;
		16'b1010101101000111: color_data = 12'b001110100111;
		16'b1010101101001000: color_data = 12'b001110100111;
		16'b1010101101001001: color_data = 12'b001110100111;
		16'b1010101101001010: color_data = 12'b001110100111;
		16'b1010101101001011: color_data = 12'b001110100111;
		16'b1010101101001100: color_data = 12'b001110100111;
		16'b1010101101001101: color_data = 12'b001110100111;
		16'b1010101101001110: color_data = 12'b001110100111;
		16'b1010101101001111: color_data = 12'b001110100111;
		16'b1010101101010000: color_data = 12'b001110100111;
		16'b1010101101010001: color_data = 12'b001110100111;
		16'b1010101101011000: color_data = 12'b001110100111;
		16'b1010101101011001: color_data = 12'b001110100111;
		16'b1010101101011010: color_data = 12'b001110100111;
		16'b1010101101011011: color_data = 12'b001110100111;
		16'b1010101101011100: color_data = 12'b001110100111;
		16'b1010101101011101: color_data = 12'b001110100111;
		16'b1010101101011110: color_data = 12'b001110100111;
		16'b1010101101011111: color_data = 12'b001110100111;
		16'b1010101101100000: color_data = 12'b001110100111;
		16'b1010101101100001: color_data = 12'b001110100111;
		16'b1010101101100010: color_data = 12'b001110100111;
		16'b1010101101100011: color_data = 12'b001110100111;
		16'b1010101101100100: color_data = 12'b001110100111;
		16'b1010101101100101: color_data = 12'b001110100111;
		16'b1010101101100110: color_data = 12'b001110100111;
		16'b1010101101100111: color_data = 12'b001110100111;
		16'b1010101101101000: color_data = 12'b001110100111;
		16'b1010101101101001: color_data = 12'b001110100111;
		16'b1010101101101010: color_data = 12'b001110100111;
		16'b1010101101101011: color_data = 12'b001110100111;
		16'b1010101101101100: color_data = 12'b001110100111;
		16'b1010101101101101: color_data = 12'b001110100111;
		16'b1010101101101110: color_data = 12'b001110100111;
		16'b1010101101101111: color_data = 12'b001110100111;
		16'b1010101101110000: color_data = 12'b001110100111;
		16'b1010101101110001: color_data = 12'b001110100111;
		16'b1010101101110010: color_data = 12'b001110100111;
		16'b1010101101110011: color_data = 12'b001110100111;
		16'b1010101101110100: color_data = 12'b001110100111;
		16'b1010101101110101: color_data = 12'b001110100111;
		16'b1010101101110110: color_data = 12'b001110100111;
		16'b1010101101110111: color_data = 12'b001110100111;
		16'b1010101101111000: color_data = 12'b001110100111;
		16'b1010101101111001: color_data = 12'b001110100111;
		16'b1010101101111010: color_data = 12'b001110100111;
		16'b1010101101111011: color_data = 12'b001110100111;
		16'b1010110000000000: color_data = 12'b001110100111;
		16'b1010110000000001: color_data = 12'b001110100111;
		16'b1010110000000010: color_data = 12'b001110100111;
		16'b1010110000000011: color_data = 12'b001110100111;
		16'b1010110000000100: color_data = 12'b001110100111;
		16'b1010110000000101: color_data = 12'b001110100111;
		16'b1010110000000110: color_data = 12'b001110100111;
		16'b1010110000000111: color_data = 12'b001110100111;
		16'b1010110000001000: color_data = 12'b001110100111;
		16'b1010110000001001: color_data = 12'b001110100111;
		16'b1010110000001010: color_data = 12'b001110100111;
		16'b1010110000001011: color_data = 12'b001110100111;
		16'b1010110000001100: color_data = 12'b001110100111;
		16'b1010110000001101: color_data = 12'b001110100111;
		16'b1010110000001110: color_data = 12'b001110100111;
		16'b1010110000001111: color_data = 12'b001110100111;
		16'b1010110000010000: color_data = 12'b001110100111;
		16'b1010110000010001: color_data = 12'b001110100111;
		16'b1010110000010010: color_data = 12'b001110100111;
		16'b1010110000010011: color_data = 12'b001110100111;
		16'b1010110000010100: color_data = 12'b001110100111;
		16'b1010110000010101: color_data = 12'b001110100111;
		16'b1010110000010110: color_data = 12'b001110100111;
		16'b1010110000010111: color_data = 12'b001110100111;
		16'b1010110000011000: color_data = 12'b001110100111;
		16'b1010110000011001: color_data = 12'b001110100111;
		16'b1010110000011010: color_data = 12'b001110100111;
		16'b1010110000011011: color_data = 12'b001110100111;
		16'b1010110000011100: color_data = 12'b001110100111;
		16'b1010110000011101: color_data = 12'b001110100111;
		16'b1010110000011110: color_data = 12'b001110100111;
		16'b1010110000011111: color_data = 12'b001110100111;
		16'b1010110000100000: color_data = 12'b001110100111;
		16'b1010110000100001: color_data = 12'b001110100111;
		16'b1010110000100010: color_data = 12'b001110100111;
		16'b1010110000100011: color_data = 12'b001110100111;
		16'b1010110000100100: color_data = 12'b001110100111;
		16'b1010110000101011: color_data = 12'b001110100111;
		16'b1010110000101100: color_data = 12'b001110100111;
		16'b1010110000101101: color_data = 12'b001110100111;
		16'b1010110000101110: color_data = 12'b001110100111;
		16'b1010110000101111: color_data = 12'b001110100111;
		16'b1010110000110000: color_data = 12'b001110100111;
		16'b1010110000110001: color_data = 12'b001110100111;
		16'b1010110000110010: color_data = 12'b001110100111;
		16'b1010110000110011: color_data = 12'b001110100111;
		16'b1010110000110100: color_data = 12'b001110100111;
		16'b1010110000110101: color_data = 12'b001110100111;
		16'b1010110000110110: color_data = 12'b001110100111;
		16'b1010110000110111: color_data = 12'b001110100111;
		16'b1010110001000100: color_data = 12'b001110100111;
		16'b1010110001000101: color_data = 12'b001110100111;
		16'b1010110001000110: color_data = 12'b001110100111;
		16'b1010110001000111: color_data = 12'b001110100111;
		16'b1010110001001000: color_data = 12'b001110100111;
		16'b1010110001001001: color_data = 12'b001110100111;
		16'b1010110001001010: color_data = 12'b001110100111;
		16'b1010110001001011: color_data = 12'b001110100111;
		16'b1010110001001100: color_data = 12'b001110100111;
		16'b1010110001001101: color_data = 12'b001110100111;
		16'b1010110001001110: color_data = 12'b001110100111;
		16'b1010110001001111: color_data = 12'b001110100111;
		16'b1010110001010110: color_data = 12'b001110100111;
		16'b1010110001010111: color_data = 12'b001110100111;
		16'b1010110001011000: color_data = 12'b001110100111;
		16'b1010110001011001: color_data = 12'b001110100111;
		16'b1010110001011010: color_data = 12'b001110100111;
		16'b1010110001011011: color_data = 12'b001110100111;
		16'b1010110001011100: color_data = 12'b001110100111;
		16'b1010110001011101: color_data = 12'b001110100111;
		16'b1010110001011110: color_data = 12'b001110100111;
		16'b1010110001011111: color_data = 12'b001110100111;
		16'b1010110001100000: color_data = 12'b001110100111;
		16'b1010110001100001: color_data = 12'b001110100111;
		16'b1010110001100010: color_data = 12'b001110100111;
		16'b1010110001100011: color_data = 12'b001110100111;
		16'b1010110001100100: color_data = 12'b001110100111;
		16'b1010110001100101: color_data = 12'b001110100111;
		16'b1010110001100110: color_data = 12'b001110100111;
		16'b1010110001100111: color_data = 12'b001110100111;
		16'b1010110001101000: color_data = 12'b001110100111;
		16'b1010110001101001: color_data = 12'b001110100111;
		16'b1010110001101010: color_data = 12'b001110100111;
		16'b1010110001101011: color_data = 12'b001110100111;
		16'b1010110001101100: color_data = 12'b001110100111;
		16'b1010110001101101: color_data = 12'b001110100111;
		16'b1010110001101110: color_data = 12'b001110100111;
		16'b1010110001110101: color_data = 12'b001110100111;
		16'b1010110001110110: color_data = 12'b001110100111;
		16'b1010110001110111: color_data = 12'b001110100111;
		16'b1010110001111000: color_data = 12'b001110100111;
		16'b1010110001111001: color_data = 12'b001110100111;
		16'b1010110001111010: color_data = 12'b001110100111;
		16'b1010110001111011: color_data = 12'b001110100111;
		16'b1010110001111100: color_data = 12'b001110100111;
		16'b1010110001111101: color_data = 12'b001110100111;
		16'b1010110001111110: color_data = 12'b001110100111;
		16'b1010110001111111: color_data = 12'b001110100111;
		16'b1010110010000000: color_data = 12'b001110100111;
		16'b1010110010001101: color_data = 12'b001110100111;
		16'b1010110010001110: color_data = 12'b001110100111;
		16'b1010110010001111: color_data = 12'b001110100111;
		16'b1010110010010000: color_data = 12'b001110100111;
		16'b1010110010010001: color_data = 12'b001110100111;
		16'b1010110010010010: color_data = 12'b001110100111;
		16'b1010110010010011: color_data = 12'b001110100111;
		16'b1010110010010100: color_data = 12'b001110100111;
		16'b1010110010010101: color_data = 12'b001110100111;
		16'b1010110010010110: color_data = 12'b001110100111;
		16'b1010110010010111: color_data = 12'b001110100111;
		16'b1010110010011000: color_data = 12'b001110100111;
		16'b1010110010011001: color_data = 12'b001110100111;
		16'b1010110010100000: color_data = 12'b001110100111;
		16'b1010110010100001: color_data = 12'b001110100111;
		16'b1010110010100010: color_data = 12'b001110100111;
		16'b1010110010100011: color_data = 12'b001110100111;
		16'b1010110010100100: color_data = 12'b001110100111;
		16'b1010110010100101: color_data = 12'b001110100111;
		16'b1010110010100110: color_data = 12'b001110100111;
		16'b1010110010100111: color_data = 12'b001110100111;
		16'b1010110010101000: color_data = 12'b001110100111;
		16'b1010110010101001: color_data = 12'b001110100111;
		16'b1010110010101010: color_data = 12'b001110100111;
		16'b1010110010101011: color_data = 12'b001110100111;
		16'b1010110010101100: color_data = 12'b001110100111;
		16'b1010110010101101: color_data = 12'b001110100111;
		16'b1010110010101110: color_data = 12'b001110100111;
		16'b1010110010101111: color_data = 12'b001110100111;
		16'b1010110010110000: color_data = 12'b001110100111;
		16'b1010110010110001: color_data = 12'b001110100111;
		16'b1010110010110010: color_data = 12'b001110100111;
		16'b1010110010110011: color_data = 12'b001110100111;
		16'b1010110010110100: color_data = 12'b001110100111;
		16'b1010110010110101: color_data = 12'b001110100111;
		16'b1010110010110110: color_data = 12'b001110100111;
		16'b1010110010110111: color_data = 12'b001110100111;
		16'b1010110010111000: color_data = 12'b001110100111;
		16'b1010110010111001: color_data = 12'b001110100111;
		16'b1010110010111010: color_data = 12'b001110100111;
		16'b1010110010111011: color_data = 12'b001110100111;
		16'b1010110010111100: color_data = 12'b001110100111;
		16'b1010110010111101: color_data = 12'b001110100111;
		16'b1010110010111110: color_data = 12'b001110100111;
		16'b1010110010111111: color_data = 12'b001110100111;
		16'b1010110011000000: color_data = 12'b001110100111;
		16'b1010110011000001: color_data = 12'b001110100111;
		16'b1010110011000010: color_data = 12'b001110100111;
		16'b1010110011000011: color_data = 12'b001110100111;
		16'b1010110011000100: color_data = 12'b001110100111;
		16'b1010110011001011: color_data = 12'b001110100111;
		16'b1010110011001100: color_data = 12'b001110100111;
		16'b1010110011001101: color_data = 12'b001110100111;
		16'b1010110011001110: color_data = 12'b001110100111;
		16'b1010110011001111: color_data = 12'b001110100111;
		16'b1010110011010000: color_data = 12'b001110100111;
		16'b1010110011010001: color_data = 12'b001110100111;
		16'b1010110011010010: color_data = 12'b001110100111;
		16'b1010110011010011: color_data = 12'b001110100111;
		16'b1010110011010100: color_data = 12'b001110100111;
		16'b1010110011010101: color_data = 12'b001110100111;
		16'b1010110011010110: color_data = 12'b001110100111;
		16'b1010110011110110: color_data = 12'b001110100111;
		16'b1010110011110111: color_data = 12'b001110100111;
		16'b1010110011111000: color_data = 12'b001110100111;
		16'b1010110011111001: color_data = 12'b001110100111;
		16'b1010110011111010: color_data = 12'b001110100111;
		16'b1010110011111011: color_data = 12'b001110100111;
		16'b1010110011111100: color_data = 12'b001110100111;
		16'b1010110011111101: color_data = 12'b001110100111;
		16'b1010110011111110: color_data = 12'b001110100111;
		16'b1010110011111111: color_data = 12'b001110100111;
		16'b1010110100000000: color_data = 12'b001110100111;
		16'b1010110100000001: color_data = 12'b001110100111;
		16'b1010110100000010: color_data = 12'b001110100111;
		16'b1010110100000011: color_data = 12'b001110100111;
		16'b1010110100000100: color_data = 12'b001110100111;
		16'b1010110100000101: color_data = 12'b001110100111;
		16'b1010110100000110: color_data = 12'b001110100111;
		16'b1010110100000111: color_data = 12'b001110100111;
		16'b1010110100001000: color_data = 12'b001110100111;
		16'b1010110100001001: color_data = 12'b001110100111;
		16'b1010110100001010: color_data = 12'b001110100111;
		16'b1010110100001011: color_data = 12'b001110100111;
		16'b1010110100001100: color_data = 12'b001110100111;
		16'b1010110100001101: color_data = 12'b001110100111;
		16'b1010110100001110: color_data = 12'b001110100111;
		16'b1010110100001111: color_data = 12'b001110100111;
		16'b1010110100010000: color_data = 12'b001110100111;
		16'b1010110100010001: color_data = 12'b001110100111;
		16'b1010110100010010: color_data = 12'b001110100111;
		16'b1010110100010011: color_data = 12'b001110100111;
		16'b1010110100010100: color_data = 12'b001110100111;
		16'b1010110100010101: color_data = 12'b001110100111;
		16'b1010110100010110: color_data = 12'b001110100111;
		16'b1010110100010111: color_data = 12'b001110100111;
		16'b1010110100011000: color_data = 12'b001110100111;
		16'b1010110100011001: color_data = 12'b001110100111;
		16'b1010110100011010: color_data = 12'b001110100111;
		16'b1010110100011011: color_data = 12'b001110100111;
		16'b1010110100011100: color_data = 12'b001110100111;
		16'b1010110100011101: color_data = 12'b001110100111;
		16'b1010110100011110: color_data = 12'b001110100111;
		16'b1010110100011111: color_data = 12'b001110100111;
		16'b1010110100100000: color_data = 12'b001110100111;
		16'b1010110100100001: color_data = 12'b001110100111;
		16'b1010110100100010: color_data = 12'b001110100111;
		16'b1010110100100011: color_data = 12'b001110100111;
		16'b1010110100100100: color_data = 12'b001110100111;
		16'b1010110100100101: color_data = 12'b001110100111;
		16'b1010110100100110: color_data = 12'b001110100111;
		16'b1010110100101101: color_data = 12'b001110100111;
		16'b1010110100101110: color_data = 12'b001110100111;
		16'b1010110100101111: color_data = 12'b001110100111;
		16'b1010110100110000: color_data = 12'b001110100111;
		16'b1010110100110001: color_data = 12'b001110100111;
		16'b1010110100110010: color_data = 12'b001110100111;
		16'b1010110100110011: color_data = 12'b001110100111;
		16'b1010110100110100: color_data = 12'b001110100111;
		16'b1010110100110101: color_data = 12'b001110100111;
		16'b1010110100110110: color_data = 12'b001110100111;
		16'b1010110100110111: color_data = 12'b001110100111;
		16'b1010110100111000: color_data = 12'b001110100111;
		16'b1010110101000101: color_data = 12'b001110100111;
		16'b1010110101000110: color_data = 12'b001110100111;
		16'b1010110101000111: color_data = 12'b001110100111;
		16'b1010110101001000: color_data = 12'b001110100111;
		16'b1010110101001001: color_data = 12'b001110100111;
		16'b1010110101001010: color_data = 12'b001110100111;
		16'b1010110101001011: color_data = 12'b001110100111;
		16'b1010110101001100: color_data = 12'b001110100111;
		16'b1010110101001101: color_data = 12'b001110100111;
		16'b1010110101001110: color_data = 12'b001110100111;
		16'b1010110101001111: color_data = 12'b001110100111;
		16'b1010110101010000: color_data = 12'b001110100111;
		16'b1010110101010001: color_data = 12'b001110100111;
		16'b1010110101011000: color_data = 12'b001110100111;
		16'b1010110101011001: color_data = 12'b001110100111;
		16'b1010110101011010: color_data = 12'b001110100111;
		16'b1010110101011011: color_data = 12'b001110100111;
		16'b1010110101011100: color_data = 12'b001110100111;
		16'b1010110101011101: color_data = 12'b001110100111;
		16'b1010110101011110: color_data = 12'b001110100111;
		16'b1010110101011111: color_data = 12'b001110100111;
		16'b1010110101100000: color_data = 12'b001110100111;
		16'b1010110101100001: color_data = 12'b001110100111;
		16'b1010110101100010: color_data = 12'b001110100111;
		16'b1010110101100011: color_data = 12'b001110100111;
		16'b1010110101100100: color_data = 12'b001110100111;
		16'b1010110101100101: color_data = 12'b001110100111;
		16'b1010110101100110: color_data = 12'b001110100111;
		16'b1010110101100111: color_data = 12'b001110100111;
		16'b1010110101101000: color_data = 12'b001110100111;
		16'b1010110101101001: color_data = 12'b001110100111;
		16'b1010110101101010: color_data = 12'b001110100111;
		16'b1010110101101011: color_data = 12'b001110100111;
		16'b1010110101101100: color_data = 12'b001110100111;
		16'b1010110101101101: color_data = 12'b001110100111;
		16'b1010110101101110: color_data = 12'b001110100111;
		16'b1010110101101111: color_data = 12'b001110100111;
		16'b1010110101110000: color_data = 12'b001110100111;
		16'b1010110101110001: color_data = 12'b001110100111;
		16'b1010110101110010: color_data = 12'b001110100111;
		16'b1010110101110011: color_data = 12'b001110100111;
		16'b1010110101110100: color_data = 12'b001110100111;
		16'b1010110101110101: color_data = 12'b001110100111;
		16'b1010110101110110: color_data = 12'b001110100111;
		16'b1010110101110111: color_data = 12'b001110100111;
		16'b1010110101111000: color_data = 12'b001110100111;
		16'b1010110101111001: color_data = 12'b001110100111;
		16'b1010110101111010: color_data = 12'b001110100111;
		16'b1010110101111011: color_data = 12'b001110100111;
		16'b1010111000000000: color_data = 12'b001110100111;
		16'b1010111000000001: color_data = 12'b001110100111;
		16'b1010111000000010: color_data = 12'b001110100111;
		16'b1010111000000011: color_data = 12'b001110100111;
		16'b1010111000000100: color_data = 12'b001110100111;
		16'b1010111000000101: color_data = 12'b001110100111;
		16'b1010111000000110: color_data = 12'b001110100111;
		16'b1010111000000111: color_data = 12'b001110100111;
		16'b1010111000001000: color_data = 12'b001110100111;
		16'b1010111000001001: color_data = 12'b001110100111;
		16'b1010111000001010: color_data = 12'b001110100111;
		16'b1010111000001011: color_data = 12'b001110100111;
		16'b1010111000001100: color_data = 12'b001110100111;
		16'b1010111000001101: color_data = 12'b001110100111;
		16'b1010111000001110: color_data = 12'b001110100111;
		16'b1010111000001111: color_data = 12'b001110100111;
		16'b1010111000010000: color_data = 12'b001110100111;
		16'b1010111000010001: color_data = 12'b001110100111;
		16'b1010111000010010: color_data = 12'b001110100111;
		16'b1010111000010011: color_data = 12'b001110100111;
		16'b1010111000010100: color_data = 12'b001110100111;
		16'b1010111000010101: color_data = 12'b001110100111;
		16'b1010111000010110: color_data = 12'b001110100111;
		16'b1010111000010111: color_data = 12'b001110100111;
		16'b1010111000011000: color_data = 12'b001110100111;
		16'b1010111000011001: color_data = 12'b001110100111;
		16'b1010111000011010: color_data = 12'b001110100111;
		16'b1010111000011011: color_data = 12'b001110100111;
		16'b1010111000011100: color_data = 12'b001110100111;
		16'b1010111000011101: color_data = 12'b001110100111;
		16'b1010111000011110: color_data = 12'b001110100111;
		16'b1010111000011111: color_data = 12'b001110100111;
		16'b1010111000100000: color_data = 12'b001110100111;
		16'b1010111000100001: color_data = 12'b001110100111;
		16'b1010111000100010: color_data = 12'b001110100111;
		16'b1010111000100011: color_data = 12'b001110100111;
		16'b1010111000100100: color_data = 12'b001110100111;
		16'b1010111000101011: color_data = 12'b001110100111;
		16'b1010111000101100: color_data = 12'b001110100111;
		16'b1010111000101101: color_data = 12'b001110100111;
		16'b1010111000101110: color_data = 12'b001110100111;
		16'b1010111000101111: color_data = 12'b001110100111;
		16'b1010111000110000: color_data = 12'b001110100111;
		16'b1010111000110001: color_data = 12'b001110100111;
		16'b1010111000110010: color_data = 12'b001110100111;
		16'b1010111000110011: color_data = 12'b001110100111;
		16'b1010111000110100: color_data = 12'b001110100111;
		16'b1010111000110101: color_data = 12'b001110100111;
		16'b1010111000110110: color_data = 12'b001110100111;
		16'b1010111000110111: color_data = 12'b001110100111;
		16'b1010111001000100: color_data = 12'b001110100111;
		16'b1010111001000101: color_data = 12'b001110100111;
		16'b1010111001000110: color_data = 12'b001110100111;
		16'b1010111001000111: color_data = 12'b001110100111;
		16'b1010111001001000: color_data = 12'b001110100111;
		16'b1010111001001001: color_data = 12'b001110100111;
		16'b1010111001001010: color_data = 12'b001110100111;
		16'b1010111001001011: color_data = 12'b001110100111;
		16'b1010111001001100: color_data = 12'b001110100111;
		16'b1010111001001101: color_data = 12'b001110100111;
		16'b1010111001001110: color_data = 12'b001110100111;
		16'b1010111001001111: color_data = 12'b001110100111;
		16'b1010111001010110: color_data = 12'b001110100111;
		16'b1010111001010111: color_data = 12'b001110100111;
		16'b1010111001011000: color_data = 12'b001110100111;
		16'b1010111001011001: color_data = 12'b001110100111;
		16'b1010111001011010: color_data = 12'b001110100111;
		16'b1010111001011011: color_data = 12'b001110100111;
		16'b1010111001011100: color_data = 12'b001110100111;
		16'b1010111001011101: color_data = 12'b001110100111;
		16'b1010111001011110: color_data = 12'b001110100111;
		16'b1010111001011111: color_data = 12'b001110100111;
		16'b1010111001100000: color_data = 12'b001110100111;
		16'b1010111001100001: color_data = 12'b001110100111;
		16'b1010111001100010: color_data = 12'b001110100111;
		16'b1010111001100011: color_data = 12'b001110100111;
		16'b1010111001100100: color_data = 12'b001110100111;
		16'b1010111001100101: color_data = 12'b001110100111;
		16'b1010111001100110: color_data = 12'b001110100111;
		16'b1010111001100111: color_data = 12'b001110100111;
		16'b1010111001101000: color_data = 12'b001110100111;
		16'b1010111001101001: color_data = 12'b001110100111;
		16'b1010111001101010: color_data = 12'b001110100111;
		16'b1010111001101011: color_data = 12'b001110100111;
		16'b1010111001101100: color_data = 12'b001110100111;
		16'b1010111001101101: color_data = 12'b001110100111;
		16'b1010111001101110: color_data = 12'b001110100111;
		16'b1010111001110101: color_data = 12'b001110100111;
		16'b1010111001110110: color_data = 12'b001110100111;
		16'b1010111001110111: color_data = 12'b001110100111;
		16'b1010111001111000: color_data = 12'b001110100111;
		16'b1010111001111001: color_data = 12'b001110100111;
		16'b1010111001111010: color_data = 12'b001110100111;
		16'b1010111001111011: color_data = 12'b001110100111;
		16'b1010111001111100: color_data = 12'b001110100111;
		16'b1010111001111101: color_data = 12'b001110100111;
		16'b1010111001111110: color_data = 12'b001110100111;
		16'b1010111001111111: color_data = 12'b001110100111;
		16'b1010111010000000: color_data = 12'b001110100111;
		16'b1010111010001101: color_data = 12'b001110100111;
		16'b1010111010001110: color_data = 12'b001110100111;
		16'b1010111010001111: color_data = 12'b001110100111;
		16'b1010111010010000: color_data = 12'b001110100111;
		16'b1010111010010001: color_data = 12'b001110100111;
		16'b1010111010010010: color_data = 12'b001110100111;
		16'b1010111010010011: color_data = 12'b001110100111;
		16'b1010111010010100: color_data = 12'b001110100111;
		16'b1010111010010101: color_data = 12'b001110100111;
		16'b1010111010010110: color_data = 12'b001110100111;
		16'b1010111010010111: color_data = 12'b001110100111;
		16'b1010111010011000: color_data = 12'b001110100111;
		16'b1010111010011001: color_data = 12'b001110100111;
		16'b1010111010100000: color_data = 12'b001110100111;
		16'b1010111010100001: color_data = 12'b001110100111;
		16'b1010111010100010: color_data = 12'b001110100111;
		16'b1010111010100011: color_data = 12'b001110100111;
		16'b1010111010100100: color_data = 12'b001110100111;
		16'b1010111010100101: color_data = 12'b001110100111;
		16'b1010111010100110: color_data = 12'b001110100111;
		16'b1010111010100111: color_data = 12'b001110100111;
		16'b1010111010101000: color_data = 12'b001110100111;
		16'b1010111010101001: color_data = 12'b001110100111;
		16'b1010111010101010: color_data = 12'b001110100111;
		16'b1010111010101011: color_data = 12'b001110100111;
		16'b1010111010101100: color_data = 12'b001110100111;
		16'b1010111010101101: color_data = 12'b001110100111;
		16'b1010111010101110: color_data = 12'b001110100111;
		16'b1010111010101111: color_data = 12'b001110100111;
		16'b1010111010110000: color_data = 12'b001110100111;
		16'b1010111010110001: color_data = 12'b001110100111;
		16'b1010111010110010: color_data = 12'b001110100111;
		16'b1010111010110011: color_data = 12'b001110100111;
		16'b1010111010110100: color_data = 12'b001110100111;
		16'b1010111010110101: color_data = 12'b001110100111;
		16'b1010111010110110: color_data = 12'b001110100111;
		16'b1010111010110111: color_data = 12'b001110100111;
		16'b1010111010111000: color_data = 12'b001110100111;
		16'b1010111010111001: color_data = 12'b001110100111;
		16'b1010111010111010: color_data = 12'b001110100111;
		16'b1010111010111011: color_data = 12'b001110100111;
		16'b1010111010111100: color_data = 12'b001110100111;
		16'b1010111010111101: color_data = 12'b001110100111;
		16'b1010111010111110: color_data = 12'b001110100111;
		16'b1010111010111111: color_data = 12'b001110100111;
		16'b1010111011000000: color_data = 12'b001110100111;
		16'b1010111011000001: color_data = 12'b001110100111;
		16'b1010111011000010: color_data = 12'b001110100111;
		16'b1010111011000011: color_data = 12'b001110100111;
		16'b1010111011000100: color_data = 12'b001110100111;
		16'b1010111011001011: color_data = 12'b001110100111;
		16'b1010111011001100: color_data = 12'b001110100111;
		16'b1010111011001101: color_data = 12'b001110100111;
		16'b1010111011001110: color_data = 12'b001110100111;
		16'b1010111011001111: color_data = 12'b001110100111;
		16'b1010111011010000: color_data = 12'b001110100111;
		16'b1010111011010001: color_data = 12'b001110100111;
		16'b1010111011010010: color_data = 12'b001110100111;
		16'b1010111011010011: color_data = 12'b001110100111;
		16'b1010111011010100: color_data = 12'b001110100111;
		16'b1010111011010101: color_data = 12'b001110100111;
		16'b1010111011010110: color_data = 12'b001110100111;
		16'b1010111011110110: color_data = 12'b001110100111;
		16'b1010111011110111: color_data = 12'b001110100111;
		16'b1010111011111000: color_data = 12'b001110100111;
		16'b1010111011111001: color_data = 12'b001110100111;
		16'b1010111011111010: color_data = 12'b001110100111;
		16'b1010111011111011: color_data = 12'b001110100111;
		16'b1010111011111100: color_data = 12'b001110100111;
		16'b1010111011111101: color_data = 12'b001110100111;
		16'b1010111011111110: color_data = 12'b001110100111;
		16'b1010111011111111: color_data = 12'b001110100111;
		16'b1010111100000000: color_data = 12'b001110100111;
		16'b1010111100000001: color_data = 12'b001110100111;
		16'b1010111100000010: color_data = 12'b001110100111;
		16'b1010111100000011: color_data = 12'b001110100111;
		16'b1010111100000100: color_data = 12'b001110100111;
		16'b1010111100000101: color_data = 12'b001110100111;
		16'b1010111100000110: color_data = 12'b001110100111;
		16'b1010111100000111: color_data = 12'b001110100111;
		16'b1010111100001000: color_data = 12'b001110100111;
		16'b1010111100001001: color_data = 12'b001110100111;
		16'b1010111100001010: color_data = 12'b001110100111;
		16'b1010111100001011: color_data = 12'b001110100111;
		16'b1010111100001100: color_data = 12'b001110100111;
		16'b1010111100001101: color_data = 12'b001110100111;
		16'b1010111100001110: color_data = 12'b001110100111;
		16'b1010111100001111: color_data = 12'b001110100111;
		16'b1010111100010000: color_data = 12'b001110100111;
		16'b1010111100010001: color_data = 12'b001110100111;
		16'b1010111100010010: color_data = 12'b001110100111;
		16'b1010111100010011: color_data = 12'b001110100111;
		16'b1010111100010100: color_data = 12'b001110100111;
		16'b1010111100010101: color_data = 12'b001110100111;
		16'b1010111100010110: color_data = 12'b001110100111;
		16'b1010111100010111: color_data = 12'b001110100111;
		16'b1010111100011000: color_data = 12'b001110100111;
		16'b1010111100011001: color_data = 12'b001110100111;
		16'b1010111100011010: color_data = 12'b001110100111;
		16'b1010111100011011: color_data = 12'b001110100111;
		16'b1010111100011100: color_data = 12'b001110100111;
		16'b1010111100011101: color_data = 12'b001110100111;
		16'b1010111100011110: color_data = 12'b001110100111;
		16'b1010111100011111: color_data = 12'b001110100111;
		16'b1010111100100000: color_data = 12'b001110100111;
		16'b1010111100100001: color_data = 12'b001110100111;
		16'b1010111100100010: color_data = 12'b001110100111;
		16'b1010111100100011: color_data = 12'b001110100111;
		16'b1010111100100100: color_data = 12'b001110100111;
		16'b1010111100100101: color_data = 12'b001110100111;
		16'b1010111100100110: color_data = 12'b001110100111;
		16'b1010111100101101: color_data = 12'b001110100111;
		16'b1010111100101110: color_data = 12'b001110100111;
		16'b1010111100101111: color_data = 12'b001110100111;
		16'b1010111100110000: color_data = 12'b001110100111;
		16'b1010111100110001: color_data = 12'b001110100111;
		16'b1010111100110010: color_data = 12'b001110100111;
		16'b1010111100110011: color_data = 12'b001110100111;
		16'b1010111100110100: color_data = 12'b001110100111;
		16'b1010111100110101: color_data = 12'b001110100111;
		16'b1010111100110110: color_data = 12'b001110100111;
		16'b1010111100110111: color_data = 12'b001110100111;
		16'b1010111100111000: color_data = 12'b001110100111;
		16'b1010111101000101: color_data = 12'b001110100111;
		16'b1010111101000110: color_data = 12'b001110100111;
		16'b1010111101000111: color_data = 12'b001110100111;
		16'b1010111101001000: color_data = 12'b001110100111;
		16'b1010111101001001: color_data = 12'b001110100111;
		16'b1010111101001010: color_data = 12'b001110100111;
		16'b1010111101001011: color_data = 12'b001110100111;
		16'b1010111101001100: color_data = 12'b001110100111;
		16'b1010111101001101: color_data = 12'b001110100111;
		16'b1010111101001110: color_data = 12'b001110100111;
		16'b1010111101001111: color_data = 12'b001110100111;
		16'b1010111101010000: color_data = 12'b001110100111;
		16'b1010111101010001: color_data = 12'b001110100111;
		16'b1010111101011000: color_data = 12'b001110100111;
		16'b1010111101011001: color_data = 12'b001110100111;
		16'b1010111101011010: color_data = 12'b001110100111;
		16'b1010111101011011: color_data = 12'b001110100111;
		16'b1010111101011100: color_data = 12'b001110100111;
		16'b1010111101011101: color_data = 12'b001110100111;
		16'b1010111101011110: color_data = 12'b001110100111;
		16'b1010111101011111: color_data = 12'b001110100111;
		16'b1010111101100000: color_data = 12'b001110100111;
		16'b1010111101100001: color_data = 12'b001110100111;
		16'b1010111101100010: color_data = 12'b001110100111;
		16'b1010111101100011: color_data = 12'b001110100111;
		16'b1010111101100100: color_data = 12'b001110100111;
		16'b1010111101100101: color_data = 12'b001110100111;
		16'b1010111101100110: color_data = 12'b001110100111;
		16'b1010111101100111: color_data = 12'b001110100111;
		16'b1010111101101000: color_data = 12'b001110100111;
		16'b1010111101101001: color_data = 12'b001110100111;
		16'b1010111101101010: color_data = 12'b001110100111;
		16'b1010111101101011: color_data = 12'b001110100111;
		16'b1010111101101100: color_data = 12'b001110100111;
		16'b1010111101101101: color_data = 12'b001110100111;
		16'b1010111101101110: color_data = 12'b001110100111;
		16'b1010111101101111: color_data = 12'b001110100111;
		16'b1010111101110000: color_data = 12'b001110100111;
		16'b1010111101110001: color_data = 12'b001110100111;
		16'b1010111101110010: color_data = 12'b001110100111;
		16'b1010111101110011: color_data = 12'b001110100111;
		16'b1010111101110100: color_data = 12'b001110100111;
		16'b1010111101110101: color_data = 12'b001110100111;
		16'b1010111101110110: color_data = 12'b001110100111;
		16'b1010111101110111: color_data = 12'b001110100111;
		16'b1010111101111000: color_data = 12'b001110100111;
		16'b1010111101111001: color_data = 12'b001110100111;
		16'b1010111101111010: color_data = 12'b001110100111;
		16'b1010111101111011: color_data = 12'b001110100111;
		16'b1011000000000000: color_data = 12'b001110100111;
		16'b1011000000000001: color_data = 12'b001110100111;
		16'b1011000000000010: color_data = 12'b001110100111;
		16'b1011000000000011: color_data = 12'b001110100111;
		16'b1011000000000100: color_data = 12'b001110100111;
		16'b1011000000000101: color_data = 12'b001110100111;
		16'b1011000000000110: color_data = 12'b001110100111;
		16'b1011000000000111: color_data = 12'b001110100111;
		16'b1011000000001000: color_data = 12'b001110100111;
		16'b1011000000001001: color_data = 12'b001110100111;
		16'b1011000000001010: color_data = 12'b001110100111;
		16'b1011000000001011: color_data = 12'b001110100111;
		16'b1011000000001100: color_data = 12'b001110100111;
		16'b1011000000001101: color_data = 12'b001110100111;
		16'b1011000000001110: color_data = 12'b001110100111;
		16'b1011000000001111: color_data = 12'b001110100111;
		16'b1011000000010000: color_data = 12'b001110100111;
		16'b1011000000010001: color_data = 12'b001110100111;
		16'b1011000000010010: color_data = 12'b001110100111;
		16'b1011000000010011: color_data = 12'b001110100111;
		16'b1011000000010100: color_data = 12'b001110100111;
		16'b1011000000010101: color_data = 12'b001110100111;
		16'b1011000000010110: color_data = 12'b001110100111;
		16'b1011000000010111: color_data = 12'b001110100111;
		16'b1011000000011000: color_data = 12'b001110100111;
		16'b1011000000011001: color_data = 12'b001110100111;
		16'b1011000000011010: color_data = 12'b001110100111;
		16'b1011000000011011: color_data = 12'b001110100111;
		16'b1011000000011100: color_data = 12'b001110100111;
		16'b1011000000011101: color_data = 12'b001110100111;
		16'b1011000000011110: color_data = 12'b001110100111;
		16'b1011000000011111: color_data = 12'b001110100111;
		16'b1011000000100000: color_data = 12'b001110100111;
		16'b1011000000100001: color_data = 12'b001110100111;
		16'b1011000000100010: color_data = 12'b001110100111;
		16'b1011000000100011: color_data = 12'b001110100111;
		16'b1011000000100100: color_data = 12'b001110100111;
		16'b1011000000101011: color_data = 12'b001110100111;
		16'b1011000000101100: color_data = 12'b001110100111;
		16'b1011000000101101: color_data = 12'b001110100111;
		16'b1011000000101110: color_data = 12'b001110100111;
		16'b1011000000101111: color_data = 12'b001110100111;
		16'b1011000000110000: color_data = 12'b001110100111;
		16'b1011000000110001: color_data = 12'b001110100111;
		16'b1011000000110010: color_data = 12'b001110100111;
		16'b1011000000110011: color_data = 12'b001110100111;
		16'b1011000000110100: color_data = 12'b001110100111;
		16'b1011000000110101: color_data = 12'b001110100111;
		16'b1011000000110110: color_data = 12'b001110100111;
		16'b1011000000110111: color_data = 12'b001110100111;
		16'b1011000001000100: color_data = 12'b001110100111;
		16'b1011000001000101: color_data = 12'b001110100111;
		16'b1011000001000110: color_data = 12'b001110100111;
		16'b1011000001000111: color_data = 12'b001110100111;
		16'b1011000001001000: color_data = 12'b001110100111;
		16'b1011000001001001: color_data = 12'b001110100111;
		16'b1011000001001010: color_data = 12'b001110100111;
		16'b1011000001001011: color_data = 12'b001110100111;
		16'b1011000001001100: color_data = 12'b001110100111;
		16'b1011000001001101: color_data = 12'b001110100111;
		16'b1011000001001110: color_data = 12'b001110100111;
		16'b1011000001001111: color_data = 12'b001110100111;
		16'b1011000001010110: color_data = 12'b001110100111;
		16'b1011000001010111: color_data = 12'b001110100111;
		16'b1011000001011000: color_data = 12'b001110100111;
		16'b1011000001011001: color_data = 12'b001110100111;
		16'b1011000001011010: color_data = 12'b001110100111;
		16'b1011000001011011: color_data = 12'b001110100111;
		16'b1011000001011100: color_data = 12'b001110100111;
		16'b1011000001011101: color_data = 12'b001110100111;
		16'b1011000001011110: color_data = 12'b001110100111;
		16'b1011000001011111: color_data = 12'b001110100111;
		16'b1011000001100000: color_data = 12'b001110100111;
		16'b1011000001100001: color_data = 12'b001110100111;
		16'b1011000001100010: color_data = 12'b001110100111;
		16'b1011000001100011: color_data = 12'b001110100111;
		16'b1011000001100100: color_data = 12'b001110100111;
		16'b1011000001100101: color_data = 12'b001110100111;
		16'b1011000001100110: color_data = 12'b001110100111;
		16'b1011000001100111: color_data = 12'b001110100111;
		16'b1011000001101000: color_data = 12'b001110100111;
		16'b1011000001101001: color_data = 12'b001110100111;
		16'b1011000001101010: color_data = 12'b001110100111;
		16'b1011000001101011: color_data = 12'b001110100111;
		16'b1011000001101100: color_data = 12'b001110100111;
		16'b1011000001101101: color_data = 12'b001110100111;
		16'b1011000001101110: color_data = 12'b001110100111;
		16'b1011000001110101: color_data = 12'b001110100111;
		16'b1011000001110110: color_data = 12'b001110100111;
		16'b1011000001110111: color_data = 12'b001110100111;
		16'b1011000001111000: color_data = 12'b001110100111;
		16'b1011000001111001: color_data = 12'b001110100111;
		16'b1011000001111010: color_data = 12'b001110100111;
		16'b1011000001111011: color_data = 12'b001110100111;
		16'b1011000001111100: color_data = 12'b001110100111;
		16'b1011000001111101: color_data = 12'b001110100111;
		16'b1011000001111110: color_data = 12'b001110100111;
		16'b1011000001111111: color_data = 12'b001110100111;
		16'b1011000010000000: color_data = 12'b001110100111;
		16'b1011000010001101: color_data = 12'b001110100111;
		16'b1011000010001110: color_data = 12'b001110100111;
		16'b1011000010001111: color_data = 12'b001110100111;
		16'b1011000010010000: color_data = 12'b001110100111;
		16'b1011000010010001: color_data = 12'b001110100111;
		16'b1011000010010010: color_data = 12'b001110100111;
		16'b1011000010010011: color_data = 12'b001110100111;
		16'b1011000010010100: color_data = 12'b001110100111;
		16'b1011000010010101: color_data = 12'b001110100111;
		16'b1011000010010110: color_data = 12'b001110100111;
		16'b1011000010010111: color_data = 12'b001110100111;
		16'b1011000010011000: color_data = 12'b001110100111;
		16'b1011000010011001: color_data = 12'b001110100111;
		16'b1011000010100000: color_data = 12'b001110100111;
		16'b1011000010100001: color_data = 12'b001110100111;
		16'b1011000010100010: color_data = 12'b001110100111;
		16'b1011000010100011: color_data = 12'b001110100111;
		16'b1011000010100100: color_data = 12'b001110100111;
		16'b1011000010100101: color_data = 12'b001110100111;
		16'b1011000010100110: color_data = 12'b001110100111;
		16'b1011000010100111: color_data = 12'b001110100111;
		16'b1011000010101000: color_data = 12'b001110100111;
		16'b1011000010101001: color_data = 12'b001110100111;
		16'b1011000010101010: color_data = 12'b001110100111;
		16'b1011000010101011: color_data = 12'b001110100111;
		16'b1011000010101100: color_data = 12'b001110100111;
		16'b1011000010101101: color_data = 12'b001110100111;
		16'b1011000010101110: color_data = 12'b001110100111;
		16'b1011000010101111: color_data = 12'b001110100111;
		16'b1011000010110000: color_data = 12'b001110100111;
		16'b1011000010110001: color_data = 12'b001110100111;
		16'b1011000010110010: color_data = 12'b001110100111;
		16'b1011000010110011: color_data = 12'b001110100111;
		16'b1011000010110100: color_data = 12'b001110100111;
		16'b1011000010110101: color_data = 12'b001110100111;
		16'b1011000010110110: color_data = 12'b001110100111;
		16'b1011000010110111: color_data = 12'b001110100111;
		16'b1011000010111000: color_data = 12'b001110100111;
		16'b1011000010111001: color_data = 12'b001110100111;
		16'b1011000010111010: color_data = 12'b001110100111;
		16'b1011000010111011: color_data = 12'b001110100111;
		16'b1011000010111100: color_data = 12'b001110100111;
		16'b1011000010111101: color_data = 12'b001110100111;
		16'b1011000010111110: color_data = 12'b001110100111;
		16'b1011000010111111: color_data = 12'b001110100111;
		16'b1011000011000000: color_data = 12'b001110100111;
		16'b1011000011000001: color_data = 12'b001110100111;
		16'b1011000011000010: color_data = 12'b001110100111;
		16'b1011000011000011: color_data = 12'b001110100111;
		16'b1011000011000100: color_data = 12'b001110100111;
		16'b1011000011001011: color_data = 12'b001110100111;
		16'b1011000011001100: color_data = 12'b001110100111;
		16'b1011000011001101: color_data = 12'b001110100111;
		16'b1011000011001110: color_data = 12'b001110100111;
		16'b1011000011001111: color_data = 12'b001110100111;
		16'b1011000011010000: color_data = 12'b001110100111;
		16'b1011000011010001: color_data = 12'b001110100111;
		16'b1011000011010010: color_data = 12'b001110100111;
		16'b1011000011010011: color_data = 12'b001110100111;
		16'b1011000011010100: color_data = 12'b001110100111;
		16'b1011000011010101: color_data = 12'b001110100111;
		16'b1011000011010110: color_data = 12'b001110100111;
		16'b1011000011110110: color_data = 12'b001110100111;
		16'b1011000011110111: color_data = 12'b001110100111;
		16'b1011000011111000: color_data = 12'b001110100111;
		16'b1011000011111001: color_data = 12'b001110100111;
		16'b1011000011111010: color_data = 12'b001110100111;
		16'b1011000011111011: color_data = 12'b001110100111;
		16'b1011000011111100: color_data = 12'b001110100111;
		16'b1011000011111101: color_data = 12'b001110100111;
		16'b1011000011111110: color_data = 12'b001110100111;
		16'b1011000011111111: color_data = 12'b001110100111;
		16'b1011000100000000: color_data = 12'b001110100111;
		16'b1011000100000001: color_data = 12'b001110100111;
		16'b1011000100000010: color_data = 12'b001110100111;
		16'b1011000100000011: color_data = 12'b001110100111;
		16'b1011000100000100: color_data = 12'b001110100111;
		16'b1011000100000101: color_data = 12'b001110100111;
		16'b1011000100000110: color_data = 12'b001110100111;
		16'b1011000100000111: color_data = 12'b001110100111;
		16'b1011000100001000: color_data = 12'b001110100111;
		16'b1011000100001001: color_data = 12'b001110100111;
		16'b1011000100001010: color_data = 12'b001110100111;
		16'b1011000100001011: color_data = 12'b001110100111;
		16'b1011000100001100: color_data = 12'b001110100111;
		16'b1011000100001101: color_data = 12'b001110100111;
		16'b1011000100001110: color_data = 12'b001110100111;
		16'b1011000100001111: color_data = 12'b001110100111;
		16'b1011000100010000: color_data = 12'b001110100111;
		16'b1011000100010001: color_data = 12'b001110100111;
		16'b1011000100010010: color_data = 12'b001110100111;
		16'b1011000100010011: color_data = 12'b001110100111;
		16'b1011000100010100: color_data = 12'b001110100111;
		16'b1011000100010101: color_data = 12'b001110100111;
		16'b1011000100010110: color_data = 12'b001110100111;
		16'b1011000100010111: color_data = 12'b001110100111;
		16'b1011000100011000: color_data = 12'b001110100111;
		16'b1011000100011001: color_data = 12'b001110100111;
		16'b1011000100011010: color_data = 12'b001110100111;
		16'b1011000100011011: color_data = 12'b001110100111;
		16'b1011000100011100: color_data = 12'b001110100111;
		16'b1011000100011101: color_data = 12'b001110100111;
		16'b1011000100011110: color_data = 12'b001110100111;
		16'b1011000100011111: color_data = 12'b001110100111;
		16'b1011000100100000: color_data = 12'b001110100111;
		16'b1011000100100001: color_data = 12'b001110100111;
		16'b1011000100100010: color_data = 12'b001110100111;
		16'b1011000100100011: color_data = 12'b001110100111;
		16'b1011000100100100: color_data = 12'b001110100111;
		16'b1011000100100101: color_data = 12'b001110100111;
		16'b1011000100100110: color_data = 12'b001110100111;
		16'b1011000100101101: color_data = 12'b001110100111;
		16'b1011000100101110: color_data = 12'b001110100111;
		16'b1011000100101111: color_data = 12'b001110100111;
		16'b1011000100110000: color_data = 12'b001110100111;
		16'b1011000100110001: color_data = 12'b001110100111;
		16'b1011000100110010: color_data = 12'b001110100111;
		16'b1011000100110011: color_data = 12'b001110100111;
		16'b1011000100110100: color_data = 12'b001110100111;
		16'b1011000100110101: color_data = 12'b001110100111;
		16'b1011000100110110: color_data = 12'b001110100111;
		16'b1011000100110111: color_data = 12'b001110100111;
		16'b1011000100111000: color_data = 12'b001110100111;
		16'b1011000101000101: color_data = 12'b001110100111;
		16'b1011000101000110: color_data = 12'b001110100111;
		16'b1011000101000111: color_data = 12'b001110100111;
		16'b1011000101001000: color_data = 12'b001110100111;
		16'b1011000101001001: color_data = 12'b001110100111;
		16'b1011000101001010: color_data = 12'b001110100111;
		16'b1011000101001011: color_data = 12'b001110100111;
		16'b1011000101001100: color_data = 12'b001110100111;
		16'b1011000101001101: color_data = 12'b001110100111;
		16'b1011000101001110: color_data = 12'b001110100111;
		16'b1011000101001111: color_data = 12'b001110100111;
		16'b1011000101010000: color_data = 12'b001110100111;
		16'b1011000101010001: color_data = 12'b001110100111;
		16'b1011000101011000: color_data = 12'b001110100111;
		16'b1011000101011001: color_data = 12'b001110100111;
		16'b1011000101011010: color_data = 12'b001110100111;
		16'b1011000101011011: color_data = 12'b001110100111;
		16'b1011000101011100: color_data = 12'b001110100111;
		16'b1011000101011101: color_data = 12'b001110100111;
		16'b1011000101011110: color_data = 12'b001110100111;
		16'b1011000101011111: color_data = 12'b001110100111;
		16'b1011000101100000: color_data = 12'b001110100111;
		16'b1011000101100001: color_data = 12'b001110100111;
		16'b1011000101100010: color_data = 12'b001110100111;
		16'b1011000101100011: color_data = 12'b001110100111;
		16'b1011000101100100: color_data = 12'b001110100111;
		16'b1011000101100101: color_data = 12'b001110100111;
		16'b1011000101100110: color_data = 12'b001110100111;
		16'b1011000101100111: color_data = 12'b001110100111;
		16'b1011000101101000: color_data = 12'b001110100111;
		16'b1011000101101001: color_data = 12'b001110100111;
		16'b1011000101101010: color_data = 12'b001110100111;
		16'b1011000101101011: color_data = 12'b001110100111;
		16'b1011000101101100: color_data = 12'b001110100111;
		16'b1011000101101101: color_data = 12'b001110100111;
		16'b1011000101101110: color_data = 12'b001110100111;
		16'b1011000101101111: color_data = 12'b001110100111;
		16'b1011000101110000: color_data = 12'b001110100111;
		16'b1011000101110001: color_data = 12'b001110100111;
		16'b1011000101110010: color_data = 12'b001110100111;
		16'b1011000101110011: color_data = 12'b001110100111;
		16'b1011000101110100: color_data = 12'b001110100111;
		16'b1011000101110101: color_data = 12'b001110100111;
		16'b1011000101110110: color_data = 12'b001110100111;
		16'b1011000101110111: color_data = 12'b001110100111;
		16'b1011000101111000: color_data = 12'b001110100111;
		16'b1011000101111001: color_data = 12'b001110100111;
		16'b1011000101111010: color_data = 12'b001110100111;
		16'b1011000101111011: color_data = 12'b001110100111;
		16'b1011001000000000: color_data = 12'b001110100111;
		16'b1011001000000001: color_data = 12'b001110100111;
		16'b1011001000000010: color_data = 12'b001110100111;
		16'b1011001000000011: color_data = 12'b001110100111;
		16'b1011001000000100: color_data = 12'b001110100111;
		16'b1011001000000101: color_data = 12'b001110100111;
		16'b1011001000000110: color_data = 12'b001110100111;
		16'b1011001000000111: color_data = 12'b001110100111;
		16'b1011001000001000: color_data = 12'b001110100111;
		16'b1011001000001001: color_data = 12'b001110100111;
		16'b1011001000001010: color_data = 12'b001110100111;
		16'b1011001000001011: color_data = 12'b001110100111;
		16'b1011001000001100: color_data = 12'b001110100111;
		16'b1011001000001101: color_data = 12'b001110100111;
		16'b1011001000001110: color_data = 12'b001110100111;
		16'b1011001000001111: color_data = 12'b001110100111;
		16'b1011001000010000: color_data = 12'b001110100111;
		16'b1011001000010001: color_data = 12'b001110100111;
		16'b1011001000010010: color_data = 12'b001110100111;
		16'b1011001000010011: color_data = 12'b001110100111;
		16'b1011001000010100: color_data = 12'b001110100111;
		16'b1011001000010101: color_data = 12'b001110100111;
		16'b1011001000010110: color_data = 12'b001110100111;
		16'b1011001000010111: color_data = 12'b001110100111;
		16'b1011001000011000: color_data = 12'b001110100111;
		16'b1011001000011001: color_data = 12'b001110100111;
		16'b1011001000011010: color_data = 12'b001110100111;
		16'b1011001000011011: color_data = 12'b001110100111;
		16'b1011001000011100: color_data = 12'b001110100111;
		16'b1011001000011101: color_data = 12'b001110100111;
		16'b1011001000011110: color_data = 12'b001110100111;
		16'b1011001000011111: color_data = 12'b001110100111;
		16'b1011001000100000: color_data = 12'b001110100111;
		16'b1011001000100001: color_data = 12'b001110100111;
		16'b1011001000100010: color_data = 12'b001110100111;
		16'b1011001000100011: color_data = 12'b001110100111;
		16'b1011001000100100: color_data = 12'b001110100111;
		16'b1011001000101011: color_data = 12'b001110100111;
		16'b1011001000101100: color_data = 12'b001110100111;
		16'b1011001000101101: color_data = 12'b001110100111;
		16'b1011001000101110: color_data = 12'b001110100111;
		16'b1011001000101111: color_data = 12'b001110100111;
		16'b1011001000110000: color_data = 12'b001110100111;
		16'b1011001000110001: color_data = 12'b001110100111;
		16'b1011001000110010: color_data = 12'b001110100111;
		16'b1011001000110011: color_data = 12'b001110100111;
		16'b1011001000110100: color_data = 12'b001110100111;
		16'b1011001000110101: color_data = 12'b001110100111;
		16'b1011001000110110: color_data = 12'b001110100111;
		16'b1011001000110111: color_data = 12'b001110100111;
		16'b1011001001000100: color_data = 12'b001110100111;
		16'b1011001001000101: color_data = 12'b001110100111;
		16'b1011001001000110: color_data = 12'b001110100111;
		16'b1011001001000111: color_data = 12'b001110100111;
		16'b1011001001001000: color_data = 12'b001110100111;
		16'b1011001001001001: color_data = 12'b001110100111;
		16'b1011001001001010: color_data = 12'b001110100111;
		16'b1011001001001011: color_data = 12'b001110100111;
		16'b1011001001001100: color_data = 12'b001110100111;
		16'b1011001001001101: color_data = 12'b001110100111;
		16'b1011001001001110: color_data = 12'b001110100111;
		16'b1011001001001111: color_data = 12'b001110100111;
		16'b1011001001010110: color_data = 12'b001110100111;
		16'b1011001001010111: color_data = 12'b001110100111;
		16'b1011001001011000: color_data = 12'b001110100111;
		16'b1011001001011001: color_data = 12'b001110100111;
		16'b1011001001011010: color_data = 12'b001110100111;
		16'b1011001001011011: color_data = 12'b001110100111;
		16'b1011001001011100: color_data = 12'b001110100111;
		16'b1011001001011101: color_data = 12'b001110100111;
		16'b1011001001011110: color_data = 12'b001110100111;
		16'b1011001001011111: color_data = 12'b001110100111;
		16'b1011001001100000: color_data = 12'b001110100111;
		16'b1011001001100001: color_data = 12'b001110100111;
		16'b1011001001100010: color_data = 12'b001110100111;
		16'b1011001001100011: color_data = 12'b001110100111;
		16'b1011001001100100: color_data = 12'b001110100111;
		16'b1011001001100101: color_data = 12'b001110100111;
		16'b1011001001100110: color_data = 12'b001110100111;
		16'b1011001001100111: color_data = 12'b001110100111;
		16'b1011001001101000: color_data = 12'b001110100111;
		16'b1011001001101001: color_data = 12'b001110100111;
		16'b1011001001101010: color_data = 12'b001110100111;
		16'b1011001001101011: color_data = 12'b001110100111;
		16'b1011001001101100: color_data = 12'b001110100111;
		16'b1011001001101101: color_data = 12'b001110100111;
		16'b1011001001101110: color_data = 12'b001110100111;
		16'b1011001001110101: color_data = 12'b001110100111;
		16'b1011001001110110: color_data = 12'b001110100111;
		16'b1011001001110111: color_data = 12'b001110100111;
		16'b1011001001111000: color_data = 12'b001110100111;
		16'b1011001001111001: color_data = 12'b001110100111;
		16'b1011001001111010: color_data = 12'b001110100111;
		16'b1011001001111011: color_data = 12'b001110100111;
		16'b1011001001111100: color_data = 12'b001110100111;
		16'b1011001001111101: color_data = 12'b001110100111;
		16'b1011001001111110: color_data = 12'b001110100111;
		16'b1011001001111111: color_data = 12'b001110100111;
		16'b1011001010000000: color_data = 12'b001110100111;
		16'b1011001010001101: color_data = 12'b001110100111;
		16'b1011001010001110: color_data = 12'b001110100111;
		16'b1011001010001111: color_data = 12'b001110100111;
		16'b1011001010010000: color_data = 12'b001110100111;
		16'b1011001010010001: color_data = 12'b001110100111;
		16'b1011001010010010: color_data = 12'b001110100111;
		16'b1011001010010011: color_data = 12'b001110100111;
		16'b1011001010010100: color_data = 12'b001110100111;
		16'b1011001010010101: color_data = 12'b001110100111;
		16'b1011001010010110: color_data = 12'b001110100111;
		16'b1011001010010111: color_data = 12'b001110100111;
		16'b1011001010011000: color_data = 12'b001110100111;
		16'b1011001010011001: color_data = 12'b001110100111;
		16'b1011001010100000: color_data = 12'b001110100111;
		16'b1011001010100001: color_data = 12'b001110100111;
		16'b1011001010100010: color_data = 12'b001110100111;
		16'b1011001010100011: color_data = 12'b001110100111;
		16'b1011001010100100: color_data = 12'b001110100111;
		16'b1011001010100101: color_data = 12'b001110100111;
		16'b1011001010100110: color_data = 12'b001110100111;
		16'b1011001010100111: color_data = 12'b001110100111;
		16'b1011001010101000: color_data = 12'b001110100111;
		16'b1011001010101001: color_data = 12'b001110100111;
		16'b1011001010101010: color_data = 12'b001110100111;
		16'b1011001010101011: color_data = 12'b001110100111;
		16'b1011001010101100: color_data = 12'b001110100111;
		16'b1011001010101101: color_data = 12'b001110100111;
		16'b1011001010101110: color_data = 12'b001110100111;
		16'b1011001010101111: color_data = 12'b001110100111;
		16'b1011001010110000: color_data = 12'b001110100111;
		16'b1011001010110001: color_data = 12'b001110100111;
		16'b1011001010110010: color_data = 12'b001110100111;
		16'b1011001010110011: color_data = 12'b001110100111;
		16'b1011001010110100: color_data = 12'b001110100111;
		16'b1011001010110101: color_data = 12'b001110100111;
		16'b1011001010110110: color_data = 12'b001110100111;
		16'b1011001010110111: color_data = 12'b001110100111;
		16'b1011001010111000: color_data = 12'b001110100111;
		16'b1011001010111001: color_data = 12'b001110100111;
		16'b1011001010111010: color_data = 12'b001110100111;
		16'b1011001010111011: color_data = 12'b001110100111;
		16'b1011001010111100: color_data = 12'b001110100111;
		16'b1011001010111101: color_data = 12'b001110100111;
		16'b1011001010111110: color_data = 12'b001110100111;
		16'b1011001010111111: color_data = 12'b001110100111;
		16'b1011001011000000: color_data = 12'b001110100111;
		16'b1011001011000001: color_data = 12'b001110100111;
		16'b1011001011000010: color_data = 12'b001110100111;
		16'b1011001011000011: color_data = 12'b001110100111;
		16'b1011001011000100: color_data = 12'b001110100111;
		16'b1011001011001011: color_data = 12'b001110100111;
		16'b1011001011001100: color_data = 12'b001110100111;
		16'b1011001011001101: color_data = 12'b001110100111;
		16'b1011001011001110: color_data = 12'b001110100111;
		16'b1011001011001111: color_data = 12'b001110100111;
		16'b1011001011010000: color_data = 12'b001110100111;
		16'b1011001011010001: color_data = 12'b001110100111;
		16'b1011001011010010: color_data = 12'b001110100111;
		16'b1011001011010011: color_data = 12'b001110100111;
		16'b1011001011010100: color_data = 12'b001110100111;
		16'b1011001011010101: color_data = 12'b001110100111;
		16'b1011001011010110: color_data = 12'b001110100111;
		16'b1011001011111100: color_data = 12'b001110100111;
		16'b1011001011111101: color_data = 12'b001110100111;
		16'b1011001011111110: color_data = 12'b001110100111;
		16'b1011001011111111: color_data = 12'b001110100111;
		16'b1011001100000000: color_data = 12'b001110100111;
		16'b1011001100000001: color_data = 12'b001110100111;
		16'b1011001100000010: color_data = 12'b001110100111;
		16'b1011001100000011: color_data = 12'b001110100111;
		16'b1011001100000100: color_data = 12'b001110100111;
		16'b1011001100000101: color_data = 12'b001110100111;
		16'b1011001100000110: color_data = 12'b001110100111;
		16'b1011001100000111: color_data = 12'b001110100111;
		16'b1011001100001000: color_data = 12'b001110100111;
		16'b1011001100001001: color_data = 12'b001110100111;
		16'b1011001100001010: color_data = 12'b001110100111;
		16'b1011001100001011: color_data = 12'b001110100111;
		16'b1011001100001100: color_data = 12'b001110100111;
		16'b1011001100001101: color_data = 12'b001110100111;
		16'b1011001100001110: color_data = 12'b001110100111;
		16'b1011001100001111: color_data = 12'b001110100111;
		16'b1011001100010000: color_data = 12'b001110100111;
		16'b1011001100010001: color_data = 12'b001110100111;
		16'b1011001100010010: color_data = 12'b001110100111;
		16'b1011001100010011: color_data = 12'b001110100111;
		16'b1011001100010100: color_data = 12'b001110100111;
		16'b1011001100010101: color_data = 12'b001110100111;
		16'b1011001100010110: color_data = 12'b001110100111;
		16'b1011001100010111: color_data = 12'b001110100111;
		16'b1011001100011000: color_data = 12'b001110100111;
		16'b1011001100011001: color_data = 12'b001110100111;
		16'b1011001100011010: color_data = 12'b001110100111;
		16'b1011001100011011: color_data = 12'b001110100111;
		16'b1011001100011100: color_data = 12'b001110100111;
		16'b1011001100011101: color_data = 12'b001110100111;
		16'b1011001100011110: color_data = 12'b001110100111;
		16'b1011001100011111: color_data = 12'b001110100111;
		16'b1011001100100000: color_data = 12'b001110100111;
		16'b1011001100101101: color_data = 12'b001110100111;
		16'b1011001100101110: color_data = 12'b001110100111;
		16'b1011001100101111: color_data = 12'b001110100111;
		16'b1011001100110000: color_data = 12'b001110100111;
		16'b1011001100110001: color_data = 12'b001110100111;
		16'b1011001100110010: color_data = 12'b001110100111;
		16'b1011001100110011: color_data = 12'b001110100111;
		16'b1011001100110100: color_data = 12'b001110100111;
		16'b1011001100110101: color_data = 12'b001110100111;
		16'b1011001100110110: color_data = 12'b001110100111;
		16'b1011001100110111: color_data = 12'b001110100111;
		16'b1011001100111000: color_data = 12'b001110100111;
		16'b1011001101000101: color_data = 12'b001110100111;
		16'b1011001101000110: color_data = 12'b001110100111;
		16'b1011001101000111: color_data = 12'b001110100111;
		16'b1011001101001000: color_data = 12'b001110100111;
		16'b1011001101001001: color_data = 12'b001110100111;
		16'b1011001101001010: color_data = 12'b001110100111;
		16'b1011001101001011: color_data = 12'b001110100111;
		16'b1011001101001100: color_data = 12'b001110100111;
		16'b1011001101001101: color_data = 12'b001110100111;
		16'b1011001101001110: color_data = 12'b001110100111;
		16'b1011001101001111: color_data = 12'b001110100111;
		16'b1011001101010000: color_data = 12'b001110100111;
		16'b1011001101010001: color_data = 12'b001110100111;
		16'b1011001101011000: color_data = 12'b001110100111;
		16'b1011001101011001: color_data = 12'b001110100111;
		16'b1011001101011010: color_data = 12'b001110100111;
		16'b1011001101011011: color_data = 12'b001110100111;
		16'b1011001101011100: color_data = 12'b001110100111;
		16'b1011001101011101: color_data = 12'b001110100111;
		16'b1011001101011110: color_data = 12'b001110100111;
		16'b1011001101011111: color_data = 12'b001110100111;
		16'b1011001101100000: color_data = 12'b001110100111;
		16'b1011001101100001: color_data = 12'b001110100111;
		16'b1011001101100010: color_data = 12'b001110100111;
		16'b1011001101100011: color_data = 12'b001110100111;
		16'b1011001101100100: color_data = 12'b001110100111;
		16'b1011001101100101: color_data = 12'b001110100111;
		16'b1011001101100110: color_data = 12'b001110100111;
		16'b1011001101100111: color_data = 12'b001110100111;
		16'b1011001101101000: color_data = 12'b001110100111;
		16'b1011001101101001: color_data = 12'b001110100111;
		16'b1011001101101010: color_data = 12'b001110100111;
		16'b1011001101101011: color_data = 12'b001110100111;
		16'b1011001101101100: color_data = 12'b001110100111;
		16'b1011001101101101: color_data = 12'b001110100111;
		16'b1011001101101110: color_data = 12'b001110100111;
		16'b1011001101101111: color_data = 12'b001110100111;
		16'b1011001101110000: color_data = 12'b001110100111;
		16'b1011001101110001: color_data = 12'b001110100111;
		16'b1011001101110010: color_data = 12'b001110100111;
		16'b1011001101110011: color_data = 12'b001110100111;
		16'b1011001101110100: color_data = 12'b001110100111;
		16'b1011001101110101: color_data = 12'b001110100111;
		16'b1011001101110110: color_data = 12'b001110100111;
		16'b1011001101110111: color_data = 12'b001110100111;
		16'b1011001101111000: color_data = 12'b001110100111;
		16'b1011001101111001: color_data = 12'b001110100111;
		16'b1011001101111010: color_data = 12'b001110100111;
		16'b1011001101111011: color_data = 12'b001110100111;
		16'b1011010000000000: color_data = 12'b001110100111;
		16'b1011010000000001: color_data = 12'b001110100111;
		16'b1011010000000010: color_data = 12'b001110100111;
		16'b1011010000000011: color_data = 12'b001110100111;
		16'b1011010000000100: color_data = 12'b001110100111;
		16'b1011010000000101: color_data = 12'b001110100111;
		16'b1011010000000110: color_data = 12'b001110100111;
		16'b1011010000000111: color_data = 12'b001110100111;
		16'b1011010000001000: color_data = 12'b001110100111;
		16'b1011010000001001: color_data = 12'b001110100111;
		16'b1011010000001010: color_data = 12'b001110100111;
		16'b1011010000001011: color_data = 12'b001110100111;
		16'b1011010000001100: color_data = 12'b001110100111;
		16'b1011010000001101: color_data = 12'b001110100111;
		16'b1011010000001110: color_data = 12'b001110100111;
		16'b1011010000001111: color_data = 12'b001110100111;
		16'b1011010000010000: color_data = 12'b001110100111;
		16'b1011010000010001: color_data = 12'b001110100111;
		16'b1011010000010010: color_data = 12'b001110100111;
		16'b1011010000010011: color_data = 12'b001110100111;
		16'b1011010000010100: color_data = 12'b001110100111;
		16'b1011010000010101: color_data = 12'b001110100111;
		16'b1011010000010110: color_data = 12'b001110100111;
		16'b1011010000010111: color_data = 12'b001110100111;
		16'b1011010000011000: color_data = 12'b001110100111;
		16'b1011010000011001: color_data = 12'b001110100111;
		16'b1011010000011010: color_data = 12'b001110100111;
		16'b1011010000011011: color_data = 12'b001110100111;
		16'b1011010000011100: color_data = 12'b001110100111;
		16'b1011010000011101: color_data = 12'b001110100111;
		16'b1011010000011110: color_data = 12'b001110100111;
		16'b1011010000011111: color_data = 12'b001110100111;
		16'b1011010000100000: color_data = 12'b001110100111;
		16'b1011010000100001: color_data = 12'b001110100111;
		16'b1011010000100010: color_data = 12'b001110100111;
		16'b1011010000100011: color_data = 12'b001110100111;
		16'b1011010000100100: color_data = 12'b001110100111;
		16'b1011010000101011: color_data = 12'b001110100111;
		16'b1011010000101100: color_data = 12'b001110100111;
		16'b1011010000101101: color_data = 12'b001110100111;
		16'b1011010000101110: color_data = 12'b001110100111;
		16'b1011010000101111: color_data = 12'b001110100111;
		16'b1011010000110000: color_data = 12'b001110100111;
		16'b1011010000110001: color_data = 12'b001110100111;
		16'b1011010000110010: color_data = 12'b001110100111;
		16'b1011010000110011: color_data = 12'b001110100111;
		16'b1011010000110100: color_data = 12'b001110100111;
		16'b1011010000110101: color_data = 12'b001110100111;
		16'b1011010000110110: color_data = 12'b001110100111;
		16'b1011010000110111: color_data = 12'b001110100111;
		16'b1011010001000100: color_data = 12'b001110100111;
		16'b1011010001000101: color_data = 12'b001110100111;
		16'b1011010001000110: color_data = 12'b001110100111;
		16'b1011010001000111: color_data = 12'b001110100111;
		16'b1011010001001000: color_data = 12'b001110100111;
		16'b1011010001001001: color_data = 12'b001110100111;
		16'b1011010001001010: color_data = 12'b001110100111;
		16'b1011010001001011: color_data = 12'b001110100111;
		16'b1011010001001100: color_data = 12'b001110100111;
		16'b1011010001001101: color_data = 12'b001110100111;
		16'b1011010001001110: color_data = 12'b001110100111;
		16'b1011010001001111: color_data = 12'b001110100111;
		16'b1011010001010110: color_data = 12'b001110100111;
		16'b1011010001010111: color_data = 12'b001110100111;
		16'b1011010001011000: color_data = 12'b001110100111;
		16'b1011010001011001: color_data = 12'b001110100111;
		16'b1011010001011010: color_data = 12'b001110100111;
		16'b1011010001011011: color_data = 12'b001110100111;
		16'b1011010001011100: color_data = 12'b001110100111;
		16'b1011010001011101: color_data = 12'b001110100111;
		16'b1011010001011110: color_data = 12'b001110100111;
		16'b1011010001011111: color_data = 12'b001110100111;
		16'b1011010001100000: color_data = 12'b001110100111;
		16'b1011010001100001: color_data = 12'b001110100111;
		16'b1011010001100010: color_data = 12'b001110100111;
		16'b1011010001100011: color_data = 12'b001110100111;
		16'b1011010001100100: color_data = 12'b001110100111;
		16'b1011010001100101: color_data = 12'b001110100111;
		16'b1011010001100110: color_data = 12'b001110100111;
		16'b1011010001100111: color_data = 12'b001110100111;
		16'b1011010001101000: color_data = 12'b001110100111;
		16'b1011010001101001: color_data = 12'b001110100111;
		16'b1011010001101010: color_data = 12'b001110100111;
		16'b1011010001101011: color_data = 12'b001110100111;
		16'b1011010001101100: color_data = 12'b001110100111;
		16'b1011010001101101: color_data = 12'b001110100111;
		16'b1011010001101110: color_data = 12'b001110100111;
		16'b1011010001110101: color_data = 12'b001110100111;
		16'b1011010001110110: color_data = 12'b001110100111;
		16'b1011010001110111: color_data = 12'b001110100111;
		16'b1011010001111000: color_data = 12'b001110100111;
		16'b1011010001111001: color_data = 12'b001110100111;
		16'b1011010001111010: color_data = 12'b001110100111;
		16'b1011010001111011: color_data = 12'b001110100111;
		16'b1011010001111100: color_data = 12'b001110100111;
		16'b1011010001111101: color_data = 12'b001110100111;
		16'b1011010001111110: color_data = 12'b001110100111;
		16'b1011010001111111: color_data = 12'b001110100111;
		16'b1011010010000000: color_data = 12'b001110100111;
		16'b1011010010001101: color_data = 12'b001110100111;
		16'b1011010010001110: color_data = 12'b001110100111;
		16'b1011010010001111: color_data = 12'b001110100111;
		16'b1011010010010000: color_data = 12'b001110100111;
		16'b1011010010010001: color_data = 12'b001110100111;
		16'b1011010010010010: color_data = 12'b001110100111;
		16'b1011010010010011: color_data = 12'b001110100111;
		16'b1011010010010100: color_data = 12'b001110100111;
		16'b1011010010010101: color_data = 12'b001110100111;
		16'b1011010010010110: color_data = 12'b001110100111;
		16'b1011010010010111: color_data = 12'b001110100111;
		16'b1011010010011000: color_data = 12'b001110100111;
		16'b1011010010011001: color_data = 12'b001110100111;
		16'b1011010010100000: color_data = 12'b001110100111;
		16'b1011010010100001: color_data = 12'b001110100111;
		16'b1011010010100010: color_data = 12'b001110100111;
		16'b1011010010100011: color_data = 12'b001110100111;
		16'b1011010010100100: color_data = 12'b001110100111;
		16'b1011010010100101: color_data = 12'b001110100111;
		16'b1011010010100110: color_data = 12'b001110100111;
		16'b1011010010100111: color_data = 12'b001110100111;
		16'b1011010010101000: color_data = 12'b001110100111;
		16'b1011010010101001: color_data = 12'b001110100111;
		16'b1011010010101010: color_data = 12'b001110100111;
		16'b1011010010101011: color_data = 12'b001110100111;
		16'b1011010010101100: color_data = 12'b001110100111;
		16'b1011010010101101: color_data = 12'b001110100111;
		16'b1011010010101110: color_data = 12'b001110100111;
		16'b1011010010101111: color_data = 12'b001110100111;
		16'b1011010010110000: color_data = 12'b001110100111;
		16'b1011010010110001: color_data = 12'b001110100111;
		16'b1011010010110010: color_data = 12'b001110100111;
		16'b1011010010110011: color_data = 12'b001110100111;
		16'b1011010010110100: color_data = 12'b001110100111;
		16'b1011010010110101: color_data = 12'b001110100111;
		16'b1011010010110110: color_data = 12'b001110100111;
		16'b1011010010110111: color_data = 12'b001110100111;
		16'b1011010010111000: color_data = 12'b001110100111;
		16'b1011010010111001: color_data = 12'b001110100111;
		16'b1011010010111010: color_data = 12'b001110100111;
		16'b1011010010111011: color_data = 12'b001110100111;
		16'b1011010010111100: color_data = 12'b001110100111;
		16'b1011010010111101: color_data = 12'b001110100111;
		16'b1011010010111110: color_data = 12'b001110100111;
		16'b1011010010111111: color_data = 12'b001110100111;
		16'b1011010011000000: color_data = 12'b001110100111;
		16'b1011010011000001: color_data = 12'b001110100111;
		16'b1011010011000010: color_data = 12'b001110100111;
		16'b1011010011000011: color_data = 12'b001110100111;
		16'b1011010011000100: color_data = 12'b001110100111;
		16'b1011010011001011: color_data = 12'b001110100111;
		16'b1011010011001100: color_data = 12'b001110100111;
		16'b1011010011001101: color_data = 12'b001110100111;
		16'b1011010011001110: color_data = 12'b001110100111;
		16'b1011010011001111: color_data = 12'b001110100111;
		16'b1011010011010000: color_data = 12'b001110100111;
		16'b1011010011010001: color_data = 12'b001110100111;
		16'b1011010011010010: color_data = 12'b001110100111;
		16'b1011010011010011: color_data = 12'b001110100111;
		16'b1011010011010100: color_data = 12'b001110100111;
		16'b1011010011010101: color_data = 12'b001110100111;
		16'b1011010011010110: color_data = 12'b001110100111;
		16'b1011010011111100: color_data = 12'b001110100111;
		16'b1011010011111101: color_data = 12'b001110100111;
		16'b1011010011111110: color_data = 12'b001110100111;
		16'b1011010011111111: color_data = 12'b001110100111;
		16'b1011010100000000: color_data = 12'b001110100111;
		16'b1011010100000001: color_data = 12'b001110100111;
		16'b1011010100000010: color_data = 12'b001110100111;
		16'b1011010100000011: color_data = 12'b001110100111;
		16'b1011010100000100: color_data = 12'b001110100111;
		16'b1011010100000101: color_data = 12'b001110100111;
		16'b1011010100000110: color_data = 12'b001110100111;
		16'b1011010100000111: color_data = 12'b001110100111;
		16'b1011010100001000: color_data = 12'b001110100111;
		16'b1011010100001001: color_data = 12'b001110100111;
		16'b1011010100001010: color_data = 12'b001110100111;
		16'b1011010100001011: color_data = 12'b001110100111;
		16'b1011010100001100: color_data = 12'b001110100111;
		16'b1011010100001101: color_data = 12'b001110100111;
		16'b1011010100001110: color_data = 12'b001110100111;
		16'b1011010100001111: color_data = 12'b001110100111;
		16'b1011010100010000: color_data = 12'b001110100111;
		16'b1011010100010001: color_data = 12'b001110100111;
		16'b1011010100010010: color_data = 12'b001110100111;
		16'b1011010100010011: color_data = 12'b001110100111;
		16'b1011010100010100: color_data = 12'b001110100111;
		16'b1011010100010101: color_data = 12'b001110100111;
		16'b1011010100010110: color_data = 12'b001110100111;
		16'b1011010100010111: color_data = 12'b001110100111;
		16'b1011010100011000: color_data = 12'b001110100111;
		16'b1011010100011001: color_data = 12'b001110100111;
		16'b1011010100011010: color_data = 12'b001110100111;
		16'b1011010100011011: color_data = 12'b001110100111;
		16'b1011010100011100: color_data = 12'b001110100111;
		16'b1011010100011101: color_data = 12'b001110100111;
		16'b1011010100011110: color_data = 12'b001110100111;
		16'b1011010100011111: color_data = 12'b001110100111;
		16'b1011010100100000: color_data = 12'b001110100111;
		16'b1011010100101101: color_data = 12'b001110100111;
		16'b1011010100101110: color_data = 12'b001110100111;
		16'b1011010100101111: color_data = 12'b001110100111;
		16'b1011010100110000: color_data = 12'b001110100111;
		16'b1011010100110001: color_data = 12'b001110100111;
		16'b1011010100110010: color_data = 12'b001110100111;
		16'b1011010100110011: color_data = 12'b001110100111;
		16'b1011010100110100: color_data = 12'b001110100111;
		16'b1011010100110101: color_data = 12'b001110100111;
		16'b1011010100110110: color_data = 12'b001110100111;
		16'b1011010100110111: color_data = 12'b001110100111;
		16'b1011010100111000: color_data = 12'b001110100111;
		16'b1011010101000101: color_data = 12'b001110100111;
		16'b1011010101000110: color_data = 12'b001110100111;
		16'b1011010101000111: color_data = 12'b001110100111;
		16'b1011010101001000: color_data = 12'b001110100111;
		16'b1011010101001001: color_data = 12'b001110100111;
		16'b1011010101001010: color_data = 12'b001110100111;
		16'b1011010101001011: color_data = 12'b001110100111;
		16'b1011010101001100: color_data = 12'b001110100111;
		16'b1011010101001101: color_data = 12'b001110100111;
		16'b1011010101001110: color_data = 12'b001110100111;
		16'b1011010101001111: color_data = 12'b001110100111;
		16'b1011010101010000: color_data = 12'b001110100111;
		16'b1011010101010001: color_data = 12'b001110100111;
		16'b1011010101011000: color_data = 12'b001110100111;
		16'b1011010101011001: color_data = 12'b001110100111;
		16'b1011010101011010: color_data = 12'b001110100111;
		16'b1011010101011011: color_data = 12'b001110100111;
		16'b1011010101011100: color_data = 12'b001110100111;
		16'b1011010101011101: color_data = 12'b001110100111;
		16'b1011010101011110: color_data = 12'b001110100111;
		16'b1011010101011111: color_data = 12'b001110100111;
		16'b1011010101100000: color_data = 12'b001110100111;
		16'b1011010101100001: color_data = 12'b001110100111;
		16'b1011010101100010: color_data = 12'b001110100111;
		16'b1011010101100011: color_data = 12'b001110100111;
		16'b1011010101100100: color_data = 12'b001110100111;
		16'b1011010101100101: color_data = 12'b001110100111;
		16'b1011010101100110: color_data = 12'b001110100111;
		16'b1011010101100111: color_data = 12'b001110100111;
		16'b1011010101101000: color_data = 12'b001110100111;
		16'b1011010101101001: color_data = 12'b001110100111;
		16'b1011010101101010: color_data = 12'b001110100111;
		16'b1011010101101011: color_data = 12'b001110100111;
		16'b1011010101101100: color_data = 12'b001110100111;
		16'b1011010101101101: color_data = 12'b001110100111;
		16'b1011010101101110: color_data = 12'b001110100111;
		16'b1011010101101111: color_data = 12'b001110100111;
		16'b1011010101110000: color_data = 12'b001110100111;
		16'b1011010101110001: color_data = 12'b001110100111;
		16'b1011010101110010: color_data = 12'b001110100111;
		16'b1011010101110011: color_data = 12'b001110100111;
		16'b1011010101110100: color_data = 12'b001110100111;
		16'b1011010101110101: color_data = 12'b001110100111;
		16'b1011010101110110: color_data = 12'b001110100111;
		16'b1011010101110111: color_data = 12'b001110100111;
		16'b1011010101111000: color_data = 12'b001110100111;
		16'b1011010101111001: color_data = 12'b001110100111;
		16'b1011010101111010: color_data = 12'b001110100111;
		16'b1011010101111011: color_data = 12'b001110100111;
		16'b1011011000000000: color_data = 12'b001110100111;
		16'b1011011000000001: color_data = 12'b001110100111;
		16'b1011011000000010: color_data = 12'b001110100111;
		16'b1011011000000011: color_data = 12'b001110100111;
		16'b1011011000000100: color_data = 12'b001110100111;
		16'b1011011000000101: color_data = 12'b001110100111;
		16'b1011011000000110: color_data = 12'b001110100111;
		16'b1011011000000111: color_data = 12'b001110100111;
		16'b1011011000001000: color_data = 12'b001110100111;
		16'b1011011000001001: color_data = 12'b001110100111;
		16'b1011011000001010: color_data = 12'b001110100111;
		16'b1011011000001011: color_data = 12'b001110100111;
		16'b1011011000001100: color_data = 12'b001110100111;
		16'b1011011000001101: color_data = 12'b001110100111;
		16'b1011011000001110: color_data = 12'b001110100111;
		16'b1011011000001111: color_data = 12'b001110100111;
		16'b1011011000010000: color_data = 12'b001110100111;
		16'b1011011000010001: color_data = 12'b001110100111;
		16'b1011011000010010: color_data = 12'b001110100111;
		16'b1011011000010011: color_data = 12'b001110100111;
		16'b1011011000010100: color_data = 12'b001110100111;
		16'b1011011000010101: color_data = 12'b001110100111;
		16'b1011011000010110: color_data = 12'b001110100111;
		16'b1011011000010111: color_data = 12'b001110100111;
		16'b1011011000011000: color_data = 12'b001110100111;
		16'b1011011000011001: color_data = 12'b001110100111;
		16'b1011011000011010: color_data = 12'b001110100111;
		16'b1011011000011011: color_data = 12'b001110100111;
		16'b1011011000011100: color_data = 12'b001110100111;
		16'b1011011000011101: color_data = 12'b001110100111;
		16'b1011011000011110: color_data = 12'b001110100111;
		16'b1011011000011111: color_data = 12'b001110100111;
		16'b1011011000100000: color_data = 12'b001110100111;
		16'b1011011000100001: color_data = 12'b001110100111;
		16'b1011011000100010: color_data = 12'b001110100111;
		16'b1011011000100011: color_data = 12'b001110100111;
		16'b1011011000100100: color_data = 12'b001110100111;
		16'b1011011000101011: color_data = 12'b001110100111;
		16'b1011011000101100: color_data = 12'b001110100111;
		16'b1011011000101101: color_data = 12'b001110100111;
		16'b1011011000101110: color_data = 12'b001110100111;
		16'b1011011000101111: color_data = 12'b001110100111;
		16'b1011011000110000: color_data = 12'b001110100111;
		16'b1011011000110001: color_data = 12'b001110100111;
		16'b1011011000110010: color_data = 12'b001110100111;
		16'b1011011000110011: color_data = 12'b001110100111;
		16'b1011011000110100: color_data = 12'b001110100111;
		16'b1011011000110101: color_data = 12'b001110100111;
		16'b1011011000110110: color_data = 12'b001110100111;
		16'b1011011000110111: color_data = 12'b001110100111;
		16'b1011011001000100: color_data = 12'b001110100111;
		16'b1011011001000101: color_data = 12'b001110100111;
		16'b1011011001000110: color_data = 12'b001110100111;
		16'b1011011001000111: color_data = 12'b001110100111;
		16'b1011011001001000: color_data = 12'b001110100111;
		16'b1011011001001001: color_data = 12'b001110100111;
		16'b1011011001001010: color_data = 12'b001110100111;
		16'b1011011001001011: color_data = 12'b001110100111;
		16'b1011011001001100: color_data = 12'b001110100111;
		16'b1011011001001101: color_data = 12'b001110100111;
		16'b1011011001001110: color_data = 12'b001110100111;
		16'b1011011001001111: color_data = 12'b001110100111;
		16'b1011011001010110: color_data = 12'b001110100111;
		16'b1011011001010111: color_data = 12'b001110100111;
		16'b1011011001011000: color_data = 12'b001110100111;
		16'b1011011001011001: color_data = 12'b001110100111;
		16'b1011011001011010: color_data = 12'b001110100111;
		16'b1011011001011011: color_data = 12'b001110100111;
		16'b1011011001011100: color_data = 12'b001110100111;
		16'b1011011001011101: color_data = 12'b001110100111;
		16'b1011011001011110: color_data = 12'b001110100111;
		16'b1011011001011111: color_data = 12'b001110100111;
		16'b1011011001100000: color_data = 12'b001110100111;
		16'b1011011001100001: color_data = 12'b001110100111;
		16'b1011011001100010: color_data = 12'b001110100111;
		16'b1011011001100011: color_data = 12'b001110100111;
		16'b1011011001100100: color_data = 12'b001110100111;
		16'b1011011001100101: color_data = 12'b001110100111;
		16'b1011011001100110: color_data = 12'b001110100111;
		16'b1011011001100111: color_data = 12'b001110100111;
		16'b1011011001101000: color_data = 12'b001110100111;
		16'b1011011001101001: color_data = 12'b001110100111;
		16'b1011011001101010: color_data = 12'b001110100111;
		16'b1011011001101011: color_data = 12'b001110100111;
		16'b1011011001101100: color_data = 12'b001110100111;
		16'b1011011001101101: color_data = 12'b001110100111;
		16'b1011011001101110: color_data = 12'b001110100111;
		16'b1011011001110101: color_data = 12'b001110100111;
		16'b1011011001110110: color_data = 12'b001110100111;
		16'b1011011001110111: color_data = 12'b001110100111;
		16'b1011011001111000: color_data = 12'b001110100111;
		16'b1011011001111001: color_data = 12'b001110100111;
		16'b1011011001111010: color_data = 12'b001110100111;
		16'b1011011001111011: color_data = 12'b001110100111;
		16'b1011011001111100: color_data = 12'b001110100111;
		16'b1011011001111101: color_data = 12'b001110100111;
		16'b1011011001111110: color_data = 12'b001110100111;
		16'b1011011001111111: color_data = 12'b001110100111;
		16'b1011011010000000: color_data = 12'b001110100111;
		16'b1011011010001101: color_data = 12'b001110100111;
		16'b1011011010001110: color_data = 12'b001110100111;
		16'b1011011010001111: color_data = 12'b001110100111;
		16'b1011011010010000: color_data = 12'b001110100111;
		16'b1011011010010001: color_data = 12'b001110100111;
		16'b1011011010010010: color_data = 12'b001110100111;
		16'b1011011010010011: color_data = 12'b001110100111;
		16'b1011011010010100: color_data = 12'b001110100111;
		16'b1011011010010101: color_data = 12'b001110100111;
		16'b1011011010010110: color_data = 12'b001110100111;
		16'b1011011010010111: color_data = 12'b001110100111;
		16'b1011011010011000: color_data = 12'b001110100111;
		16'b1011011010011001: color_data = 12'b001110100111;
		16'b1011011010100000: color_data = 12'b001110100111;
		16'b1011011010100001: color_data = 12'b001110100111;
		16'b1011011010100010: color_data = 12'b001110100111;
		16'b1011011010100011: color_data = 12'b001110100111;
		16'b1011011010100100: color_data = 12'b001110100111;
		16'b1011011010100101: color_data = 12'b001110100111;
		16'b1011011010100110: color_data = 12'b001110100111;
		16'b1011011010100111: color_data = 12'b001110100111;
		16'b1011011010101000: color_data = 12'b001110100111;
		16'b1011011010101001: color_data = 12'b001110100111;
		16'b1011011010101010: color_data = 12'b001110100111;
		16'b1011011010101011: color_data = 12'b001110100111;
		16'b1011011010101100: color_data = 12'b001110100111;
		16'b1011011010101101: color_data = 12'b001110100111;
		16'b1011011010101110: color_data = 12'b001110100111;
		16'b1011011010101111: color_data = 12'b001110100111;
		16'b1011011010110000: color_data = 12'b001110100111;
		16'b1011011010110001: color_data = 12'b001110100111;
		16'b1011011010110010: color_data = 12'b001110100111;
		16'b1011011010110011: color_data = 12'b001110100111;
		16'b1011011010110100: color_data = 12'b001110100111;
		16'b1011011010110101: color_data = 12'b001110100111;
		16'b1011011010110110: color_data = 12'b001110100111;
		16'b1011011010110111: color_data = 12'b001110100111;
		16'b1011011010111000: color_data = 12'b001110100111;
		16'b1011011010111001: color_data = 12'b001110100111;
		16'b1011011010111010: color_data = 12'b001110100111;
		16'b1011011010111011: color_data = 12'b001110100111;
		16'b1011011010111100: color_data = 12'b001110100111;
		16'b1011011010111101: color_data = 12'b001110100111;
		16'b1011011010111110: color_data = 12'b001110100111;
		16'b1011011010111111: color_data = 12'b001110100111;
		16'b1011011011000000: color_data = 12'b001110100111;
		16'b1011011011000001: color_data = 12'b001110100111;
		16'b1011011011000010: color_data = 12'b001110100111;
		16'b1011011011000011: color_data = 12'b001110100111;
		16'b1011011011000100: color_data = 12'b001110100111;
		16'b1011011011001011: color_data = 12'b001110100111;
		16'b1011011011001100: color_data = 12'b001110100111;
		16'b1011011011001101: color_data = 12'b001110100111;
		16'b1011011011001110: color_data = 12'b001110100111;
		16'b1011011011001111: color_data = 12'b001110100111;
		16'b1011011011010000: color_data = 12'b001110100111;
		16'b1011011011010001: color_data = 12'b001110100111;
		16'b1011011011010010: color_data = 12'b001110100111;
		16'b1011011011010011: color_data = 12'b001110100111;
		16'b1011011011010100: color_data = 12'b001110100111;
		16'b1011011011010101: color_data = 12'b001110100111;
		16'b1011011011010110: color_data = 12'b001110100111;
		16'b1011011011111100: color_data = 12'b001110100111;
		16'b1011011011111101: color_data = 12'b001110100111;
		16'b1011011011111110: color_data = 12'b001110100111;
		16'b1011011011111111: color_data = 12'b001110100111;
		16'b1011011100000000: color_data = 12'b001110100111;
		16'b1011011100000001: color_data = 12'b001110100111;
		16'b1011011100000010: color_data = 12'b001110100111;
		16'b1011011100000011: color_data = 12'b001110100111;
		16'b1011011100000100: color_data = 12'b001110100111;
		16'b1011011100000101: color_data = 12'b001110100111;
		16'b1011011100000110: color_data = 12'b001110100111;
		16'b1011011100000111: color_data = 12'b001110100111;
		16'b1011011100001000: color_data = 12'b001110100111;
		16'b1011011100001001: color_data = 12'b001110100111;
		16'b1011011100001010: color_data = 12'b001110100111;
		16'b1011011100001011: color_data = 12'b001110100111;
		16'b1011011100001100: color_data = 12'b001110100111;
		16'b1011011100001101: color_data = 12'b001110100111;
		16'b1011011100001110: color_data = 12'b001110100111;
		16'b1011011100001111: color_data = 12'b001110100111;
		16'b1011011100010000: color_data = 12'b001110100111;
		16'b1011011100010001: color_data = 12'b001110100111;
		16'b1011011100010010: color_data = 12'b001110100111;
		16'b1011011100010011: color_data = 12'b001110100111;
		16'b1011011100010100: color_data = 12'b001110100111;
		16'b1011011100010101: color_data = 12'b001110100111;
		16'b1011011100010110: color_data = 12'b001110100111;
		16'b1011011100010111: color_data = 12'b001110100111;
		16'b1011011100011000: color_data = 12'b001110100111;
		16'b1011011100011001: color_data = 12'b001110100111;
		16'b1011011100011010: color_data = 12'b001110100111;
		16'b1011011100011011: color_data = 12'b001110100111;
		16'b1011011100011100: color_data = 12'b001110100111;
		16'b1011011100011101: color_data = 12'b001110100111;
		16'b1011011100011110: color_data = 12'b001110100111;
		16'b1011011100011111: color_data = 12'b001110100111;
		16'b1011011100100000: color_data = 12'b001110100111;
		16'b1011011100101101: color_data = 12'b001110100111;
		16'b1011011100101110: color_data = 12'b001110100111;
		16'b1011011100101111: color_data = 12'b001110100111;
		16'b1011011100110000: color_data = 12'b001110100111;
		16'b1011011100110001: color_data = 12'b001110100111;
		16'b1011011100110010: color_data = 12'b001110100111;
		16'b1011011100110011: color_data = 12'b001110100111;
		16'b1011011100110100: color_data = 12'b001110100111;
		16'b1011011100110101: color_data = 12'b001110100111;
		16'b1011011100110110: color_data = 12'b001110100111;
		16'b1011011100110111: color_data = 12'b001110100111;
		16'b1011011100111000: color_data = 12'b001110100111;
		16'b1011011101000101: color_data = 12'b001110100111;
		16'b1011011101000110: color_data = 12'b001110100111;
		16'b1011011101000111: color_data = 12'b001110100111;
		16'b1011011101001000: color_data = 12'b001110100111;
		16'b1011011101001001: color_data = 12'b001110100111;
		16'b1011011101001010: color_data = 12'b001110100111;
		16'b1011011101001011: color_data = 12'b001110100111;
		16'b1011011101001100: color_data = 12'b001110100111;
		16'b1011011101001101: color_data = 12'b001110100111;
		16'b1011011101001110: color_data = 12'b001110100111;
		16'b1011011101001111: color_data = 12'b001110100111;
		16'b1011011101010000: color_data = 12'b001110100111;
		16'b1011011101010001: color_data = 12'b001110100111;
		16'b1011011101011000: color_data = 12'b001110100111;
		16'b1011011101011001: color_data = 12'b001110100111;
		16'b1011011101011010: color_data = 12'b001110100111;
		16'b1011011101011011: color_data = 12'b001110100111;
		16'b1011011101011100: color_data = 12'b001110100111;
		16'b1011011101011101: color_data = 12'b001110100111;
		16'b1011011101011110: color_data = 12'b001110100111;
		16'b1011011101011111: color_data = 12'b001110100111;
		16'b1011011101100000: color_data = 12'b001110100111;
		16'b1011011101100001: color_data = 12'b001110100111;
		16'b1011011101100010: color_data = 12'b001110100111;
		16'b1011011101100011: color_data = 12'b001110100111;
		16'b1011011101100100: color_data = 12'b001110100111;
		16'b1011011101100101: color_data = 12'b001110100111;
		16'b1011011101100110: color_data = 12'b001110100111;
		16'b1011011101100111: color_data = 12'b001110100111;
		16'b1011011101101000: color_data = 12'b001110100111;
		16'b1011011101101001: color_data = 12'b001110100111;
		16'b1011011101101010: color_data = 12'b001110100111;
		16'b1011011101101011: color_data = 12'b001110100111;
		16'b1011011101101100: color_data = 12'b001110100111;
		16'b1011011101101101: color_data = 12'b001110100111;
		16'b1011011101101110: color_data = 12'b001110100111;
		16'b1011011101101111: color_data = 12'b001110100111;
		16'b1011011101110000: color_data = 12'b001110100111;
		16'b1011011101110001: color_data = 12'b001110100111;
		16'b1011011101110010: color_data = 12'b001110100111;
		16'b1011011101110011: color_data = 12'b001110100111;
		16'b1011011101110100: color_data = 12'b001110100111;
		16'b1011011101110101: color_data = 12'b001110100111;
		16'b1011011101110110: color_data = 12'b001110100111;
		16'b1011011101110111: color_data = 12'b001110100111;
		16'b1011011101111000: color_data = 12'b001110100111;
		16'b1011011101111001: color_data = 12'b001110100111;
		16'b1011011101111010: color_data = 12'b001110100111;
		16'b1011011101111011: color_data = 12'b001110100111;
		16'b1011100000000000: color_data = 12'b001110100111;
		16'b1011100000000001: color_data = 12'b001110100111;
		16'b1011100000000010: color_data = 12'b001110100111;
		16'b1011100000000011: color_data = 12'b001110100111;
		16'b1011100000000100: color_data = 12'b001110100111;
		16'b1011100000000101: color_data = 12'b001110100111;
		16'b1011100000000110: color_data = 12'b001110100111;
		16'b1011100000000111: color_data = 12'b001110100111;
		16'b1011100000001000: color_data = 12'b001110100111;
		16'b1011100000001001: color_data = 12'b001110100111;
		16'b1011100000001010: color_data = 12'b001110100111;
		16'b1011100000001011: color_data = 12'b001110100111;
		16'b1011100000001100: color_data = 12'b001110100111;
		16'b1011100000001101: color_data = 12'b001110100111;
		16'b1011100000001110: color_data = 12'b001110100111;
		16'b1011100000001111: color_data = 12'b001110100111;
		16'b1011100000010000: color_data = 12'b001110100111;
		16'b1011100000010001: color_data = 12'b001110100111;
		16'b1011100000010010: color_data = 12'b001110100111;
		16'b1011100000010011: color_data = 12'b001110100111;
		16'b1011100000010100: color_data = 12'b001110100111;
		16'b1011100000010101: color_data = 12'b001110100111;
		16'b1011100000010110: color_data = 12'b001110100111;
		16'b1011100000010111: color_data = 12'b001110100111;
		16'b1011100000011000: color_data = 12'b001110100111;
		16'b1011100000011001: color_data = 12'b001110100111;
		16'b1011100000011010: color_data = 12'b001110100111;
		16'b1011100000011011: color_data = 12'b001110100111;
		16'b1011100000011100: color_data = 12'b001110100111;
		16'b1011100000011101: color_data = 12'b001110100111;
		16'b1011100000011110: color_data = 12'b001110100111;
		16'b1011100000011111: color_data = 12'b001110100111;
		16'b1011100000100000: color_data = 12'b001110100111;
		16'b1011100000100001: color_data = 12'b001110100111;
		16'b1011100000100010: color_data = 12'b001110100111;
		16'b1011100000100011: color_data = 12'b001110100111;
		16'b1011100000100100: color_data = 12'b001110100111;
		16'b1011100000101011: color_data = 12'b001110100111;
		16'b1011100000101100: color_data = 12'b001110100111;
		16'b1011100000101101: color_data = 12'b001110100111;
		16'b1011100000101110: color_data = 12'b001110100111;
		16'b1011100000101111: color_data = 12'b001110100111;
		16'b1011100000110000: color_data = 12'b001110100111;
		16'b1011100000110001: color_data = 12'b001110100111;
		16'b1011100000110010: color_data = 12'b001110100111;
		16'b1011100000110011: color_data = 12'b001110100111;
		16'b1011100000110100: color_data = 12'b001110100111;
		16'b1011100000110101: color_data = 12'b001110100111;
		16'b1011100000110110: color_data = 12'b001110100111;
		16'b1011100000110111: color_data = 12'b001110100111;
		16'b1011100001000100: color_data = 12'b001110100111;
		16'b1011100001000101: color_data = 12'b001110100111;
		16'b1011100001000110: color_data = 12'b001110100111;
		16'b1011100001000111: color_data = 12'b001110100111;
		16'b1011100001001000: color_data = 12'b001110100111;
		16'b1011100001001001: color_data = 12'b001110100111;
		16'b1011100001001010: color_data = 12'b001110100111;
		16'b1011100001001011: color_data = 12'b001110100111;
		16'b1011100001001100: color_data = 12'b001110100111;
		16'b1011100001001101: color_data = 12'b001110100111;
		16'b1011100001001110: color_data = 12'b001110100111;
		16'b1011100001001111: color_data = 12'b001110100111;
		16'b1011100001010110: color_data = 12'b001110100111;
		16'b1011100001010111: color_data = 12'b001110100111;
		16'b1011100001011000: color_data = 12'b001110100111;
		16'b1011100001011001: color_data = 12'b001110100111;
		16'b1011100001011010: color_data = 12'b001110100111;
		16'b1011100001011011: color_data = 12'b001110100111;
		16'b1011100001011100: color_data = 12'b001110100111;
		16'b1011100001011101: color_data = 12'b001110100111;
		16'b1011100001011110: color_data = 12'b001110100111;
		16'b1011100001011111: color_data = 12'b001110100111;
		16'b1011100001100000: color_data = 12'b001110100111;
		16'b1011100001100001: color_data = 12'b001110100111;
		16'b1011100001100010: color_data = 12'b001110100111;
		16'b1011100001100011: color_data = 12'b001110100111;
		16'b1011100001100100: color_data = 12'b001110100111;
		16'b1011100001100101: color_data = 12'b001110100111;
		16'b1011100001100110: color_data = 12'b001110100111;
		16'b1011100001100111: color_data = 12'b001110100111;
		16'b1011100001101000: color_data = 12'b001110100111;
		16'b1011100001101001: color_data = 12'b001110100111;
		16'b1011100001101010: color_data = 12'b001110100111;
		16'b1011100001101011: color_data = 12'b001110100111;
		16'b1011100001101100: color_data = 12'b001110100111;
		16'b1011100001101101: color_data = 12'b001110100111;
		16'b1011100001101110: color_data = 12'b001110100111;
		16'b1011100001110101: color_data = 12'b001110100111;
		16'b1011100001110110: color_data = 12'b001110100111;
		16'b1011100001110111: color_data = 12'b001110100111;
		16'b1011100001111000: color_data = 12'b001110100111;
		16'b1011100001111001: color_data = 12'b001110100111;
		16'b1011100001111010: color_data = 12'b001110100111;
		16'b1011100001111011: color_data = 12'b001110100111;
		16'b1011100001111100: color_data = 12'b001110100111;
		16'b1011100001111101: color_data = 12'b001110100111;
		16'b1011100001111110: color_data = 12'b001110100111;
		16'b1011100001111111: color_data = 12'b001110100111;
		16'b1011100010000000: color_data = 12'b001110100111;
		16'b1011100010001101: color_data = 12'b001110100111;
		16'b1011100010001110: color_data = 12'b001110100111;
		16'b1011100010001111: color_data = 12'b001110100111;
		16'b1011100010010000: color_data = 12'b001110100111;
		16'b1011100010010001: color_data = 12'b001110100111;
		16'b1011100010010010: color_data = 12'b001110100111;
		16'b1011100010010011: color_data = 12'b001110100111;
		16'b1011100010010100: color_data = 12'b001110100111;
		16'b1011100010010101: color_data = 12'b001110100111;
		16'b1011100010010110: color_data = 12'b001110100111;
		16'b1011100010010111: color_data = 12'b001110100111;
		16'b1011100010011000: color_data = 12'b001110100111;
		16'b1011100010011001: color_data = 12'b001110100111;
		16'b1011100010100000: color_data = 12'b001110100111;
		16'b1011100010100001: color_data = 12'b001110100111;
		16'b1011100010100010: color_data = 12'b001110100111;
		16'b1011100010100011: color_data = 12'b001110100111;
		16'b1011100010100100: color_data = 12'b001110100111;
		16'b1011100010100101: color_data = 12'b001110100111;
		16'b1011100010100110: color_data = 12'b001110100111;
		16'b1011100010100111: color_data = 12'b001110100111;
		16'b1011100010101000: color_data = 12'b001110100111;
		16'b1011100010101001: color_data = 12'b001110100111;
		16'b1011100010101010: color_data = 12'b001110100111;
		16'b1011100010101011: color_data = 12'b001110100111;
		16'b1011100010101100: color_data = 12'b001110100111;
		16'b1011100010101101: color_data = 12'b001110100111;
		16'b1011100010101110: color_data = 12'b001110100111;
		16'b1011100010101111: color_data = 12'b001110100111;
		16'b1011100010110000: color_data = 12'b001110100111;
		16'b1011100010110001: color_data = 12'b001110100111;
		16'b1011100010110010: color_data = 12'b001110100111;
		16'b1011100010110011: color_data = 12'b001110100111;
		16'b1011100010110100: color_data = 12'b001110100111;
		16'b1011100010110101: color_data = 12'b001110100111;
		16'b1011100010110110: color_data = 12'b001110100111;
		16'b1011100010110111: color_data = 12'b001110100111;
		16'b1011100010111000: color_data = 12'b001110100111;
		16'b1011100010111001: color_data = 12'b001110100111;
		16'b1011100010111010: color_data = 12'b001110100111;
		16'b1011100010111011: color_data = 12'b001110100111;
		16'b1011100010111100: color_data = 12'b001110100111;
		16'b1011100010111101: color_data = 12'b001110100111;
		16'b1011100010111110: color_data = 12'b001110100111;
		16'b1011100010111111: color_data = 12'b001110100111;
		16'b1011100011000000: color_data = 12'b001110100111;
		16'b1011100011000001: color_data = 12'b001110100111;
		16'b1011100011000010: color_data = 12'b001110100111;
		16'b1011100011000011: color_data = 12'b001110100111;
		16'b1011100011000100: color_data = 12'b001110100111;
		16'b1011100011001011: color_data = 12'b001110100111;
		16'b1011100011001100: color_data = 12'b001110100111;
		16'b1011100011001101: color_data = 12'b001110100111;
		16'b1011100011001110: color_data = 12'b001110100111;
		16'b1011100011001111: color_data = 12'b001110100111;
		16'b1011100011010000: color_data = 12'b001110100111;
		16'b1011100011010001: color_data = 12'b001110100111;
		16'b1011100011010010: color_data = 12'b001110100111;
		16'b1011100011010011: color_data = 12'b001110100111;
		16'b1011100011010100: color_data = 12'b001110100111;
		16'b1011100011010101: color_data = 12'b001110100111;
		16'b1011100011010110: color_data = 12'b001110100111;
		16'b1011100011111100: color_data = 12'b001110100111;
		16'b1011100011111101: color_data = 12'b001110100111;
		16'b1011100011111110: color_data = 12'b001110100111;
		16'b1011100011111111: color_data = 12'b001110100111;
		16'b1011100100000000: color_data = 12'b001110100111;
		16'b1011100100000001: color_data = 12'b001110100111;
		16'b1011100100000010: color_data = 12'b001110100111;
		16'b1011100100000011: color_data = 12'b001110100111;
		16'b1011100100000100: color_data = 12'b001110100111;
		16'b1011100100000101: color_data = 12'b001110100111;
		16'b1011100100000110: color_data = 12'b001110100111;
		16'b1011100100000111: color_data = 12'b001110100111;
		16'b1011100100001000: color_data = 12'b001110100111;
		16'b1011100100001001: color_data = 12'b001110100111;
		16'b1011100100001010: color_data = 12'b001110100111;
		16'b1011100100001011: color_data = 12'b001110100111;
		16'b1011100100001100: color_data = 12'b001110100111;
		16'b1011100100001101: color_data = 12'b001110100111;
		16'b1011100100001110: color_data = 12'b001110100111;
		16'b1011100100001111: color_data = 12'b001110100111;
		16'b1011100100010000: color_data = 12'b001110100111;
		16'b1011100100010001: color_data = 12'b001110100111;
		16'b1011100100010010: color_data = 12'b001110100111;
		16'b1011100100010011: color_data = 12'b001110100111;
		16'b1011100100010100: color_data = 12'b001110100111;
		16'b1011100100010101: color_data = 12'b001110100111;
		16'b1011100100010110: color_data = 12'b001110100111;
		16'b1011100100010111: color_data = 12'b001110100111;
		16'b1011100100011000: color_data = 12'b001110100111;
		16'b1011100100011001: color_data = 12'b001110100111;
		16'b1011100100011010: color_data = 12'b001110100111;
		16'b1011100100011011: color_data = 12'b001110100111;
		16'b1011100100011100: color_data = 12'b001110100111;
		16'b1011100100011101: color_data = 12'b001110100111;
		16'b1011100100011110: color_data = 12'b001110100111;
		16'b1011100100011111: color_data = 12'b001110100111;
		16'b1011100100100000: color_data = 12'b001110100111;
		16'b1011100100101101: color_data = 12'b001110100111;
		16'b1011100100101110: color_data = 12'b001110100111;
		16'b1011100100101111: color_data = 12'b001110100111;
		16'b1011100100110000: color_data = 12'b001110100111;
		16'b1011100100110001: color_data = 12'b001110100111;
		16'b1011100100110010: color_data = 12'b001110100111;
		16'b1011100100110011: color_data = 12'b001110100111;
		16'b1011100100110100: color_data = 12'b001110100111;
		16'b1011100100110101: color_data = 12'b001110100111;
		16'b1011100100110110: color_data = 12'b001110100111;
		16'b1011100100110111: color_data = 12'b001110100111;
		16'b1011100100111000: color_data = 12'b001110100111;
		16'b1011100101000101: color_data = 12'b001110100111;
		16'b1011100101000110: color_data = 12'b001110100111;
		16'b1011100101000111: color_data = 12'b001110100111;
		16'b1011100101001000: color_data = 12'b001110100111;
		16'b1011100101001001: color_data = 12'b001110100111;
		16'b1011100101001010: color_data = 12'b001110100111;
		16'b1011100101001011: color_data = 12'b001110100111;
		16'b1011100101001100: color_data = 12'b001110100111;
		16'b1011100101001101: color_data = 12'b001110100111;
		16'b1011100101001110: color_data = 12'b001110100111;
		16'b1011100101001111: color_data = 12'b001110100111;
		16'b1011100101010000: color_data = 12'b001110100111;
		16'b1011100101010001: color_data = 12'b001110100111;
		16'b1011100101011000: color_data = 12'b001110100111;
		16'b1011100101011001: color_data = 12'b001110100111;
		16'b1011100101011010: color_data = 12'b001110100111;
		16'b1011100101011011: color_data = 12'b001110100111;
		16'b1011100101011100: color_data = 12'b001110100111;
		16'b1011100101011101: color_data = 12'b001110100111;
		16'b1011100101011110: color_data = 12'b001110100111;
		16'b1011100101011111: color_data = 12'b001110100111;
		16'b1011100101100000: color_data = 12'b001110100111;
		16'b1011100101100001: color_data = 12'b001110100111;
		16'b1011100101100010: color_data = 12'b001110100111;
		16'b1011100101100011: color_data = 12'b001110100111;
		16'b1011100101100100: color_data = 12'b001110100111;
		16'b1011100101100101: color_data = 12'b001110100111;
		16'b1011100101100110: color_data = 12'b001110100111;
		16'b1011100101100111: color_data = 12'b001110100111;
		16'b1011100101101000: color_data = 12'b001110100111;
		16'b1011100101101001: color_data = 12'b001110100111;
		16'b1011100101101010: color_data = 12'b001110100111;
		16'b1011100101101011: color_data = 12'b001110100111;
		16'b1011100101101100: color_data = 12'b001110100111;
		16'b1011100101101101: color_data = 12'b001110100111;
		16'b1011100101101110: color_data = 12'b001110100111;
		16'b1011100101101111: color_data = 12'b001110100111;
		16'b1011100101110000: color_data = 12'b001110100111;
		16'b1011100101110001: color_data = 12'b001110100111;
		16'b1011100101110010: color_data = 12'b001110100111;
		16'b1011100101110011: color_data = 12'b001110100111;
		16'b1011100101110100: color_data = 12'b001110100111;
		16'b1011100101110101: color_data = 12'b001110100111;
		16'b1011100101110110: color_data = 12'b001110100111;
		16'b1011100101110111: color_data = 12'b001110100111;
		16'b1011100101111000: color_data = 12'b001110100111;
		16'b1011100101111001: color_data = 12'b001110100111;
		16'b1011100101111010: color_data = 12'b001110100111;
		16'b1011100101111011: color_data = 12'b001110100111;
		16'b1011101000000000: color_data = 12'b001110100111;
		16'b1011101000000001: color_data = 12'b001110100111;
		16'b1011101000000010: color_data = 12'b001110100111;
		16'b1011101000000011: color_data = 12'b001110100111;
		16'b1011101000000100: color_data = 12'b001110100111;
		16'b1011101000000101: color_data = 12'b001110100111;
		16'b1011101000000110: color_data = 12'b001110100111;
		16'b1011101000000111: color_data = 12'b001110100111;
		16'b1011101000001000: color_data = 12'b001110100111;
		16'b1011101000001001: color_data = 12'b001110100111;
		16'b1011101000001010: color_data = 12'b001110100111;
		16'b1011101000001011: color_data = 12'b001110100111;
		16'b1011101000001100: color_data = 12'b001110100111;
		16'b1011101000001101: color_data = 12'b001110100111;
		16'b1011101000001110: color_data = 12'b001110100111;
		16'b1011101000001111: color_data = 12'b001110100111;
		16'b1011101000010000: color_data = 12'b001110100111;
		16'b1011101000010001: color_data = 12'b001110100111;
		16'b1011101000010010: color_data = 12'b001110100111;
		16'b1011101000010011: color_data = 12'b001110100111;
		16'b1011101000010100: color_data = 12'b001110100111;
		16'b1011101000010101: color_data = 12'b001110100111;
		16'b1011101000010110: color_data = 12'b001110100111;
		16'b1011101000010111: color_data = 12'b001110100111;
		16'b1011101000011000: color_data = 12'b001110100111;
		16'b1011101000011001: color_data = 12'b001110100111;
		16'b1011101000011010: color_data = 12'b001110100111;
		16'b1011101000011011: color_data = 12'b001110100111;
		16'b1011101000011100: color_data = 12'b001110100111;
		16'b1011101000011101: color_data = 12'b001110100111;
		16'b1011101000011110: color_data = 12'b001110100111;
		16'b1011101000011111: color_data = 12'b001110100111;
		16'b1011101000100000: color_data = 12'b001110100111;
		16'b1011101000100001: color_data = 12'b001110100111;
		16'b1011101000100010: color_data = 12'b001110100111;
		16'b1011101000100011: color_data = 12'b001110100111;
		16'b1011101000100100: color_data = 12'b001110100111;
		16'b1011101000101011: color_data = 12'b001110100111;
		16'b1011101000101100: color_data = 12'b001110100111;
		16'b1011101000101101: color_data = 12'b001110100111;
		16'b1011101000101110: color_data = 12'b001110100111;
		16'b1011101000101111: color_data = 12'b001110100111;
		16'b1011101000110000: color_data = 12'b001110100111;
		16'b1011101000110001: color_data = 12'b001110100111;
		16'b1011101000110010: color_data = 12'b001110100111;
		16'b1011101000110011: color_data = 12'b001110100111;
		16'b1011101000110100: color_data = 12'b001110100111;
		16'b1011101000110101: color_data = 12'b001110100111;
		16'b1011101000110110: color_data = 12'b001110100111;
		16'b1011101000110111: color_data = 12'b001110100111;
		16'b1011101001000100: color_data = 12'b001110100111;
		16'b1011101001000101: color_data = 12'b001110100111;
		16'b1011101001000110: color_data = 12'b001110100111;
		16'b1011101001000111: color_data = 12'b001110100111;
		16'b1011101001001000: color_data = 12'b001110100111;
		16'b1011101001001001: color_data = 12'b001110100111;
		16'b1011101001001010: color_data = 12'b001110100111;
		16'b1011101001001011: color_data = 12'b001110100111;
		16'b1011101001001100: color_data = 12'b001110100111;
		16'b1011101001001101: color_data = 12'b001110100111;
		16'b1011101001001110: color_data = 12'b001110100111;
		16'b1011101001001111: color_data = 12'b001110100111;
		16'b1011101001010110: color_data = 12'b001110100111;
		16'b1011101001010111: color_data = 12'b001110100111;
		16'b1011101001011000: color_data = 12'b001110100111;
		16'b1011101001011001: color_data = 12'b001110100111;
		16'b1011101001011010: color_data = 12'b001110100111;
		16'b1011101001011011: color_data = 12'b001110100111;
		16'b1011101001011100: color_data = 12'b001110100111;
		16'b1011101001011101: color_data = 12'b001110100111;
		16'b1011101001011110: color_data = 12'b001110100111;
		16'b1011101001011111: color_data = 12'b001110100111;
		16'b1011101001100000: color_data = 12'b001110100111;
		16'b1011101001100001: color_data = 12'b001110100111;
		16'b1011101001100010: color_data = 12'b001110100111;
		16'b1011101001100011: color_data = 12'b001110100111;
		16'b1011101001100100: color_data = 12'b001110100111;
		16'b1011101001100101: color_data = 12'b001110100111;
		16'b1011101001100110: color_data = 12'b001110100111;
		16'b1011101001100111: color_data = 12'b001110100111;
		16'b1011101001101000: color_data = 12'b001110100111;
		16'b1011101001101001: color_data = 12'b001110100111;
		16'b1011101001101010: color_data = 12'b001110100111;
		16'b1011101001101011: color_data = 12'b001110100111;
		16'b1011101001101100: color_data = 12'b001110100111;
		16'b1011101001101101: color_data = 12'b001110100111;
		16'b1011101001101110: color_data = 12'b001110100111;
		16'b1011101001110101: color_data = 12'b001110100111;
		16'b1011101001110110: color_data = 12'b001110100111;
		16'b1011101001110111: color_data = 12'b001110100111;
		16'b1011101001111000: color_data = 12'b001110100111;
		16'b1011101001111001: color_data = 12'b001110100111;
		16'b1011101001111010: color_data = 12'b001110100111;
		16'b1011101001111011: color_data = 12'b001110100111;
		16'b1011101001111100: color_data = 12'b001110100111;
		16'b1011101001111101: color_data = 12'b001110100111;
		16'b1011101001111110: color_data = 12'b001110100111;
		16'b1011101001111111: color_data = 12'b001110100111;
		16'b1011101010000000: color_data = 12'b001110100111;
		16'b1011101010001101: color_data = 12'b001110100111;
		16'b1011101010001110: color_data = 12'b001110100111;
		16'b1011101010001111: color_data = 12'b001110100111;
		16'b1011101010010000: color_data = 12'b001110100111;
		16'b1011101010010001: color_data = 12'b001110100111;
		16'b1011101010010010: color_data = 12'b001110100111;
		16'b1011101010010011: color_data = 12'b001110100111;
		16'b1011101010010100: color_data = 12'b001110100111;
		16'b1011101010010101: color_data = 12'b001110100111;
		16'b1011101010010110: color_data = 12'b001110100111;
		16'b1011101010010111: color_data = 12'b001110100111;
		16'b1011101010011000: color_data = 12'b001110100111;
		16'b1011101010011001: color_data = 12'b001110100111;
		16'b1011101010100000: color_data = 12'b001110100111;
		16'b1011101010100001: color_data = 12'b001110100111;
		16'b1011101010100010: color_data = 12'b001110100111;
		16'b1011101010100011: color_data = 12'b001110100111;
		16'b1011101010100100: color_data = 12'b001110100111;
		16'b1011101010100101: color_data = 12'b001110100111;
		16'b1011101010100110: color_data = 12'b001110100111;
		16'b1011101010100111: color_data = 12'b001110100111;
		16'b1011101010101000: color_data = 12'b001110100111;
		16'b1011101010101001: color_data = 12'b001110100111;
		16'b1011101010101010: color_data = 12'b001110100111;
		16'b1011101010101011: color_data = 12'b001110100111;
		16'b1011101010101100: color_data = 12'b001110100111;
		16'b1011101010101101: color_data = 12'b001110100111;
		16'b1011101010101110: color_data = 12'b001110100111;
		16'b1011101010101111: color_data = 12'b001110100111;
		16'b1011101010110000: color_data = 12'b001110100111;
		16'b1011101010110001: color_data = 12'b001110100111;
		16'b1011101010110010: color_data = 12'b001110100111;
		16'b1011101010110011: color_data = 12'b001110100111;
		16'b1011101010110100: color_data = 12'b001110100111;
		16'b1011101010110101: color_data = 12'b001110100111;
		16'b1011101010110110: color_data = 12'b001110100111;
		16'b1011101010110111: color_data = 12'b001110100111;
		16'b1011101010111000: color_data = 12'b001110100111;
		16'b1011101010111001: color_data = 12'b001110100111;
		16'b1011101010111010: color_data = 12'b001110100111;
		16'b1011101010111011: color_data = 12'b001110100111;
		16'b1011101010111100: color_data = 12'b001110100111;
		16'b1011101010111101: color_data = 12'b001110100111;
		16'b1011101010111110: color_data = 12'b001110100111;
		16'b1011101010111111: color_data = 12'b001110100111;
		16'b1011101011000000: color_data = 12'b001110100111;
		16'b1011101011000001: color_data = 12'b001110100111;
		16'b1011101011000010: color_data = 12'b001110100111;
		16'b1011101011000011: color_data = 12'b001110100111;
		16'b1011101011000100: color_data = 12'b001110100111;
		16'b1011101011001011: color_data = 12'b001110100111;
		16'b1011101011001100: color_data = 12'b001110100111;
		16'b1011101011001101: color_data = 12'b001110100111;
		16'b1011101011001110: color_data = 12'b001110100111;
		16'b1011101011001111: color_data = 12'b001110100111;
		16'b1011101011010000: color_data = 12'b001110100111;
		16'b1011101011010001: color_data = 12'b001110100111;
		16'b1011101011010010: color_data = 12'b001110100111;
		16'b1011101011010011: color_data = 12'b001110100111;
		16'b1011101011010100: color_data = 12'b001110100111;
		16'b1011101011010101: color_data = 12'b001110100111;
		16'b1011101011010110: color_data = 12'b001110100111;
		16'b1011101011111100: color_data = 12'b001110100111;
		16'b1011101011111101: color_data = 12'b001110100111;
		16'b1011101011111110: color_data = 12'b001110100111;
		16'b1011101011111111: color_data = 12'b001110100111;
		16'b1011101100000000: color_data = 12'b001110100111;
		16'b1011101100000001: color_data = 12'b001110100111;
		16'b1011101100000010: color_data = 12'b001110100111;
		16'b1011101100000011: color_data = 12'b001110100111;
		16'b1011101100000100: color_data = 12'b001110100111;
		16'b1011101100000101: color_data = 12'b001110100111;
		16'b1011101100000110: color_data = 12'b001110100111;
		16'b1011101100000111: color_data = 12'b001110100111;
		16'b1011101100001000: color_data = 12'b001110100111;
		16'b1011101100001001: color_data = 12'b001110100111;
		16'b1011101100001010: color_data = 12'b001110100111;
		16'b1011101100001011: color_data = 12'b001110100111;
		16'b1011101100001100: color_data = 12'b001110100111;
		16'b1011101100001101: color_data = 12'b001110100111;
		16'b1011101100001110: color_data = 12'b001110100111;
		16'b1011101100001111: color_data = 12'b001110100111;
		16'b1011101100010000: color_data = 12'b001110100111;
		16'b1011101100010001: color_data = 12'b001110100111;
		16'b1011101100010010: color_data = 12'b001110100111;
		16'b1011101100010011: color_data = 12'b001110100111;
		16'b1011101100010100: color_data = 12'b001110100111;
		16'b1011101100010101: color_data = 12'b001110100111;
		16'b1011101100010110: color_data = 12'b001110100111;
		16'b1011101100010111: color_data = 12'b001110100111;
		16'b1011101100011000: color_data = 12'b001110100111;
		16'b1011101100011001: color_data = 12'b001110100111;
		16'b1011101100011010: color_data = 12'b001110100111;
		16'b1011101100011011: color_data = 12'b001110100111;
		16'b1011101100011100: color_data = 12'b001110100111;
		16'b1011101100011101: color_data = 12'b001110100111;
		16'b1011101100011110: color_data = 12'b001110100111;
		16'b1011101100011111: color_data = 12'b001110100111;
		16'b1011101100100000: color_data = 12'b001110100111;
		16'b1011101100101101: color_data = 12'b001110100111;
		16'b1011101100101110: color_data = 12'b001110100111;
		16'b1011101100101111: color_data = 12'b001110100111;
		16'b1011101100110000: color_data = 12'b001110100111;
		16'b1011101100110001: color_data = 12'b001110100111;
		16'b1011101100110010: color_data = 12'b001110100111;
		16'b1011101100110011: color_data = 12'b001110100111;
		16'b1011101100110100: color_data = 12'b001110100111;
		16'b1011101100110101: color_data = 12'b001110100111;
		16'b1011101100110110: color_data = 12'b001110100111;
		16'b1011101100110111: color_data = 12'b001110100111;
		16'b1011101100111000: color_data = 12'b001110100111;
		16'b1011101101000101: color_data = 12'b001110100111;
		16'b1011101101000110: color_data = 12'b001110100111;
		16'b1011101101000111: color_data = 12'b001110100111;
		16'b1011101101001000: color_data = 12'b001110100111;
		16'b1011101101001001: color_data = 12'b001110100111;
		16'b1011101101001010: color_data = 12'b001110100111;
		16'b1011101101001011: color_data = 12'b001110100111;
		16'b1011101101001100: color_data = 12'b001110100111;
		16'b1011101101001101: color_data = 12'b001110100111;
		16'b1011101101001110: color_data = 12'b001110100111;
		16'b1011101101001111: color_data = 12'b001110100111;
		16'b1011101101010000: color_data = 12'b001110100111;
		16'b1011101101010001: color_data = 12'b001110100111;
		16'b1011101101011000: color_data = 12'b001110100111;
		16'b1011101101011001: color_data = 12'b001110100111;
		16'b1011101101011010: color_data = 12'b001110100111;
		16'b1011101101011011: color_data = 12'b001110100111;
		16'b1011101101011100: color_data = 12'b001110100111;
		16'b1011101101011101: color_data = 12'b001110100111;
		16'b1011101101011110: color_data = 12'b001110100111;
		16'b1011101101011111: color_data = 12'b001110100111;
		16'b1011101101100000: color_data = 12'b001110100111;
		16'b1011101101100001: color_data = 12'b001110100111;
		16'b1011101101100010: color_data = 12'b001110100111;
		16'b1011101101100011: color_data = 12'b001110100111;
		16'b1011101101100100: color_data = 12'b001110100111;
		16'b1011101101100101: color_data = 12'b001110100111;
		16'b1011101101100110: color_data = 12'b001110100111;
		16'b1011101101100111: color_data = 12'b001110100111;
		16'b1011101101101000: color_data = 12'b001110100111;
		16'b1011101101101001: color_data = 12'b001110100111;
		16'b1011101101101010: color_data = 12'b001110100111;
		16'b1011101101101011: color_data = 12'b001110100111;
		16'b1011101101101100: color_data = 12'b001110100111;
		16'b1011101101101101: color_data = 12'b001110100111;
		16'b1011101101101110: color_data = 12'b001110100111;
		16'b1011101101101111: color_data = 12'b001110100111;
		16'b1011101101110000: color_data = 12'b001110100111;
		16'b1011101101110001: color_data = 12'b001110100111;
		16'b1011101101110010: color_data = 12'b001110100111;
		16'b1011101101110011: color_data = 12'b001110100111;
		16'b1011101101110100: color_data = 12'b001110100111;
		16'b1011101101110101: color_data = 12'b001110100111;
		16'b1011101101110110: color_data = 12'b001110100111;
		16'b1011101101110111: color_data = 12'b001110100111;
		16'b1011101101111000: color_data = 12'b001110100111;
		16'b1011101101111001: color_data = 12'b001110100111;
		16'b1011101101111010: color_data = 12'b001110100111;
		16'b1011101101111011: color_data = 12'b001110100111;
		16'b1011110000000000: color_data = 12'b001110100111;
		16'b1011110000000001: color_data = 12'b001110100111;
		16'b1011110000000010: color_data = 12'b001110100111;
		16'b1011110000000011: color_data = 12'b001110100111;
		16'b1011110000000100: color_data = 12'b001110100111;
		16'b1011110000000101: color_data = 12'b001110100111;
		16'b1011110000000110: color_data = 12'b001110100111;
		16'b1011110000000111: color_data = 12'b001110100111;
		16'b1011110000001000: color_data = 12'b001110100111;
		16'b1011110000001001: color_data = 12'b001110100111;
		16'b1011110000001010: color_data = 12'b001110100111;
		16'b1011110000001011: color_data = 12'b001110100111;
		16'b1011110000001100: color_data = 12'b001110100111;
		16'b1011110000001101: color_data = 12'b001110100111;
		16'b1011110000001110: color_data = 12'b001110100111;
		16'b1011110000001111: color_data = 12'b001110100111;
		16'b1011110000010000: color_data = 12'b001110100111;
		16'b1011110000010001: color_data = 12'b001110100111;
		16'b1011110000010010: color_data = 12'b001110100111;
		16'b1011110000010011: color_data = 12'b001110100111;
		16'b1011110000010100: color_data = 12'b001110100111;
		16'b1011110000010101: color_data = 12'b001110100111;
		16'b1011110000010110: color_data = 12'b001110100111;
		16'b1011110000010111: color_data = 12'b001110100111;
		16'b1011110000011000: color_data = 12'b001110100111;
		16'b1011110000011001: color_data = 12'b001110100111;
		16'b1011110000011010: color_data = 12'b001110100111;
		16'b1011110000011011: color_data = 12'b001110100111;
		16'b1011110000011100: color_data = 12'b001110100111;
		16'b1011110000011101: color_data = 12'b001110100111;
		16'b1011110000011110: color_data = 12'b001110100111;
		16'b1011110000011111: color_data = 12'b001110100111;
		16'b1011110000100000: color_data = 12'b001110100111;
		16'b1011110000100001: color_data = 12'b001110100111;
		16'b1011110000100010: color_data = 12'b001110100111;
		16'b1011110000100011: color_data = 12'b001110100111;
		16'b1011110000100100: color_data = 12'b001110100111;
		16'b1011110000101011: color_data = 12'b001110100111;
		16'b1011110000101100: color_data = 12'b001110100111;
		16'b1011110000101101: color_data = 12'b001110100111;
		16'b1011110000101110: color_data = 12'b001110100111;
		16'b1011110000101111: color_data = 12'b001110100111;
		16'b1011110000110000: color_data = 12'b001110100111;
		16'b1011110000110001: color_data = 12'b001110100111;
		16'b1011110000110010: color_data = 12'b001110100111;
		16'b1011110000110011: color_data = 12'b001110100111;
		16'b1011110000110100: color_data = 12'b001110100111;
		16'b1011110000110101: color_data = 12'b001110100111;
		16'b1011110000110110: color_data = 12'b001110100111;
		16'b1011110000110111: color_data = 12'b001110100111;
		16'b1011110001000100: color_data = 12'b001110100111;
		16'b1011110001000101: color_data = 12'b001110100111;
		16'b1011110001000110: color_data = 12'b001110100111;
		16'b1011110001000111: color_data = 12'b001110100111;
		16'b1011110001001000: color_data = 12'b001110100111;
		16'b1011110001001001: color_data = 12'b001110100111;
		16'b1011110001001010: color_data = 12'b001110100111;
		16'b1011110001001011: color_data = 12'b001110100111;
		16'b1011110001001100: color_data = 12'b001110100111;
		16'b1011110001001101: color_data = 12'b001110100111;
		16'b1011110001001110: color_data = 12'b001110100111;
		16'b1011110001001111: color_data = 12'b001110100111;
		16'b1011110001010110: color_data = 12'b001110100111;
		16'b1011110001010111: color_data = 12'b001110100111;
		16'b1011110001011000: color_data = 12'b001110100111;
		16'b1011110001011001: color_data = 12'b001110100111;
		16'b1011110001011010: color_data = 12'b001110100111;
		16'b1011110001011011: color_data = 12'b001110100111;
		16'b1011110001011100: color_data = 12'b001110100111;
		16'b1011110001011101: color_data = 12'b001110100111;
		16'b1011110001011110: color_data = 12'b001110100111;
		16'b1011110001011111: color_data = 12'b001110100111;
		16'b1011110001100000: color_data = 12'b001110100111;
		16'b1011110001100001: color_data = 12'b001110100111;
		16'b1011110001100010: color_data = 12'b001110100111;
		16'b1011110001100011: color_data = 12'b001110100111;
		16'b1011110001100100: color_data = 12'b001110100111;
		16'b1011110001100101: color_data = 12'b001110100111;
		16'b1011110001100110: color_data = 12'b001110100111;
		16'b1011110001100111: color_data = 12'b001110100111;
		16'b1011110001101000: color_data = 12'b001110100111;
		16'b1011110001101001: color_data = 12'b001110100111;
		16'b1011110001101010: color_data = 12'b001110100111;
		16'b1011110001101011: color_data = 12'b001110100111;
		16'b1011110001101100: color_data = 12'b001110100111;
		16'b1011110001101101: color_data = 12'b001110100111;
		16'b1011110001101110: color_data = 12'b001110100111;
		16'b1011110001110101: color_data = 12'b001110100111;
		16'b1011110001110110: color_data = 12'b001110100111;
		16'b1011110001110111: color_data = 12'b001110100111;
		16'b1011110001111000: color_data = 12'b001110100111;
		16'b1011110001111001: color_data = 12'b001110100111;
		16'b1011110001111010: color_data = 12'b001110100111;
		16'b1011110001111011: color_data = 12'b001110100111;
		16'b1011110001111100: color_data = 12'b001110100111;
		16'b1011110001111101: color_data = 12'b001110100111;
		16'b1011110001111110: color_data = 12'b001110100111;
		16'b1011110001111111: color_data = 12'b001110100111;
		16'b1011110010000000: color_data = 12'b001110100111;
		16'b1011110010001101: color_data = 12'b001110100111;
		16'b1011110010001110: color_data = 12'b001110100111;
		16'b1011110010001111: color_data = 12'b001110100111;
		16'b1011110010010000: color_data = 12'b001110100111;
		16'b1011110010010001: color_data = 12'b001110100111;
		16'b1011110010010010: color_data = 12'b001110100111;
		16'b1011110010010011: color_data = 12'b001110100111;
		16'b1011110010010100: color_data = 12'b001110100111;
		16'b1011110010010101: color_data = 12'b001110100111;
		16'b1011110010010110: color_data = 12'b001110100111;
		16'b1011110010010111: color_data = 12'b001110100111;
		16'b1011110010011000: color_data = 12'b001110100111;
		16'b1011110010011001: color_data = 12'b001110100111;
		16'b1011110010100000: color_data = 12'b001110100111;
		16'b1011110010100001: color_data = 12'b001110100111;
		16'b1011110010100010: color_data = 12'b001110100111;
		16'b1011110010100011: color_data = 12'b001110100111;
		16'b1011110010100100: color_data = 12'b001110100111;
		16'b1011110010100101: color_data = 12'b001110100111;
		16'b1011110010100110: color_data = 12'b001110100111;
		16'b1011110010100111: color_data = 12'b001110100111;
		16'b1011110010101000: color_data = 12'b001110100111;
		16'b1011110010101001: color_data = 12'b001110100111;
		16'b1011110010101010: color_data = 12'b001110100111;
		16'b1011110010101011: color_data = 12'b001110100111;
		16'b1011110010101100: color_data = 12'b001110100111;
		16'b1011110010101101: color_data = 12'b001110100111;
		16'b1011110010101110: color_data = 12'b001110100111;
		16'b1011110010101111: color_data = 12'b001110100111;
		16'b1011110010110000: color_data = 12'b001110100111;
		16'b1011110010110001: color_data = 12'b001110100111;
		16'b1011110010110010: color_data = 12'b001110100111;
		16'b1011110010110011: color_data = 12'b001110100111;
		16'b1011110010110100: color_data = 12'b001110100111;
		16'b1011110010110101: color_data = 12'b001110100111;
		16'b1011110010110110: color_data = 12'b001110100111;
		16'b1011110010110111: color_data = 12'b001110100111;
		16'b1011110010111000: color_data = 12'b001110100111;
		16'b1011110010111001: color_data = 12'b001110100111;
		16'b1011110010111010: color_data = 12'b001110100111;
		16'b1011110010111011: color_data = 12'b001110100111;
		16'b1011110010111100: color_data = 12'b001110100111;
		16'b1011110010111101: color_data = 12'b001110100111;
		16'b1011110010111110: color_data = 12'b001110100111;
		16'b1011110010111111: color_data = 12'b001110100111;
		16'b1011110011000000: color_data = 12'b001110100111;
		16'b1011110011000001: color_data = 12'b001110100111;
		16'b1011110011000010: color_data = 12'b001110100111;
		16'b1011110011000011: color_data = 12'b001110100111;
		16'b1011110011000100: color_data = 12'b001110100111;
		16'b1011110011001011: color_data = 12'b001110100111;
		16'b1011110011001100: color_data = 12'b001110100111;
		16'b1011110011001101: color_data = 12'b001110100111;
		16'b1011110011001110: color_data = 12'b001110100111;
		16'b1011110011001111: color_data = 12'b001110100111;
		16'b1011110011010000: color_data = 12'b001110100111;
		16'b1011110011010001: color_data = 12'b001110100111;
		16'b1011110011010010: color_data = 12'b001110100111;
		16'b1011110011010011: color_data = 12'b001110100111;
		16'b1011110011010100: color_data = 12'b001110100111;
		16'b1011110011010101: color_data = 12'b001110100111;
		16'b1011110011010110: color_data = 12'b001110100111;
		16'b1011110011111100: color_data = 12'b001110100111;
		16'b1011110011111101: color_data = 12'b001110100111;
		16'b1011110011111110: color_data = 12'b001110100111;
		16'b1011110011111111: color_data = 12'b001110100111;
		16'b1011110100000000: color_data = 12'b001110100111;
		16'b1011110100000001: color_data = 12'b001110100111;
		16'b1011110100000010: color_data = 12'b001110100111;
		16'b1011110100000011: color_data = 12'b001110100111;
		16'b1011110100000100: color_data = 12'b001110100111;
		16'b1011110100000101: color_data = 12'b001110100111;
		16'b1011110100000110: color_data = 12'b001110100111;
		16'b1011110100000111: color_data = 12'b001110100111;
		16'b1011110100001000: color_data = 12'b001110100111;
		16'b1011110100001001: color_data = 12'b001110100111;
		16'b1011110100001010: color_data = 12'b001110100111;
		16'b1011110100001011: color_data = 12'b001110100111;
		16'b1011110100001100: color_data = 12'b001110100111;
		16'b1011110100001101: color_data = 12'b001110100111;
		16'b1011110100001110: color_data = 12'b001110100111;
		16'b1011110100001111: color_data = 12'b001110100111;
		16'b1011110100010000: color_data = 12'b001110100111;
		16'b1011110100010001: color_data = 12'b001110100111;
		16'b1011110100010010: color_data = 12'b001110100111;
		16'b1011110100010011: color_data = 12'b001110100111;
		16'b1011110100010100: color_data = 12'b001110100111;
		16'b1011110100010101: color_data = 12'b001110100111;
		16'b1011110100010110: color_data = 12'b001110100111;
		16'b1011110100010111: color_data = 12'b001110100111;
		16'b1011110100011000: color_data = 12'b001110100111;
		16'b1011110100011001: color_data = 12'b001110100111;
		16'b1011110100011010: color_data = 12'b001110100111;
		16'b1011110100011011: color_data = 12'b001110100111;
		16'b1011110100011100: color_data = 12'b001110100111;
		16'b1011110100011101: color_data = 12'b001110100111;
		16'b1011110100011110: color_data = 12'b001110100111;
		16'b1011110100011111: color_data = 12'b001110100111;
		16'b1011110100100000: color_data = 12'b001110100111;
		16'b1011110100101101: color_data = 12'b001110100111;
		16'b1011110100101110: color_data = 12'b001110100111;
		16'b1011110100101111: color_data = 12'b001110100111;
		16'b1011110100110000: color_data = 12'b001110100111;
		16'b1011110100110001: color_data = 12'b001110100111;
		16'b1011110100110010: color_data = 12'b001110100111;
		16'b1011110100110011: color_data = 12'b001110100111;
		16'b1011110100110100: color_data = 12'b001110100111;
		16'b1011110100110101: color_data = 12'b001110100111;
		16'b1011110100110110: color_data = 12'b001110100111;
		16'b1011110100110111: color_data = 12'b001110100111;
		16'b1011110100111000: color_data = 12'b001110100111;
		16'b1011110101000101: color_data = 12'b001110100111;
		16'b1011110101000110: color_data = 12'b001110100111;
		16'b1011110101000111: color_data = 12'b001110100111;
		16'b1011110101001000: color_data = 12'b001110100111;
		16'b1011110101001001: color_data = 12'b001110100111;
		16'b1011110101001010: color_data = 12'b001110100111;
		16'b1011110101001011: color_data = 12'b001110100111;
		16'b1011110101001100: color_data = 12'b001110100111;
		16'b1011110101001101: color_data = 12'b001110100111;
		16'b1011110101001110: color_data = 12'b001110100111;
		16'b1011110101001111: color_data = 12'b001110100111;
		16'b1011110101010000: color_data = 12'b001110100111;
		16'b1011110101010001: color_data = 12'b001110100111;
		16'b1011110101011000: color_data = 12'b001110100111;
		16'b1011110101011001: color_data = 12'b001110100111;
		16'b1011110101011010: color_data = 12'b001110100111;
		16'b1011110101011011: color_data = 12'b001110100111;
		16'b1011110101011100: color_data = 12'b001110100111;
		16'b1011110101011101: color_data = 12'b001110100111;
		16'b1011110101011110: color_data = 12'b001110100111;
		16'b1011110101011111: color_data = 12'b001110100111;
		16'b1011110101100000: color_data = 12'b001110100111;
		16'b1011110101100001: color_data = 12'b001110100111;
		16'b1011110101100010: color_data = 12'b001110100111;
		16'b1011110101100011: color_data = 12'b001110100111;
		16'b1011110101100100: color_data = 12'b001110100111;
		16'b1011110101100101: color_data = 12'b001110100111;
		16'b1011110101100110: color_data = 12'b001110100111;
		16'b1011110101100111: color_data = 12'b001110100111;
		16'b1011110101101000: color_data = 12'b001110100111;
		16'b1011110101101001: color_data = 12'b001110100111;
		16'b1011110101101010: color_data = 12'b001110100111;
		16'b1011110101101011: color_data = 12'b001110100111;
		16'b1011110101101100: color_data = 12'b001110100111;
		16'b1011110101101101: color_data = 12'b001110100111;
		16'b1011110101101110: color_data = 12'b001110100111;
		16'b1011110101101111: color_data = 12'b001110100111;
		16'b1011110101110000: color_data = 12'b001110100111;
		16'b1011110101110001: color_data = 12'b001110100111;
		16'b1011110101110010: color_data = 12'b001110100111;
		16'b1011110101110011: color_data = 12'b001110100111;
		16'b1011110101110100: color_data = 12'b001110100111;
		16'b1011110101110101: color_data = 12'b001110100111;
		16'b1011110101110110: color_data = 12'b001110100111;
		16'b1011110101110111: color_data = 12'b001110100111;
		16'b1011110101111000: color_data = 12'b001110100111;
		16'b1011110101111001: color_data = 12'b001110100111;
		16'b1011110101111010: color_data = 12'b001110100111;
		16'b1011110101111011: color_data = 12'b001110100111;
		16'b1011111000000000: color_data = 12'b001110100111;
		16'b1011111000000001: color_data = 12'b001110100111;
		16'b1011111000000010: color_data = 12'b001110100111;
		16'b1011111000000011: color_data = 12'b001110100111;
		16'b1011111000000100: color_data = 12'b001110100111;
		16'b1011111000000101: color_data = 12'b001110100111;
		16'b1011111000000110: color_data = 12'b001110100111;
		16'b1011111000000111: color_data = 12'b001110100111;
		16'b1011111000001000: color_data = 12'b001110100111;
		16'b1011111000001001: color_data = 12'b001110100111;
		16'b1011111000001010: color_data = 12'b001110100111;
		16'b1011111000001011: color_data = 12'b001110100111;
		16'b1011111000001100: color_data = 12'b001110100111;
		16'b1011111000001101: color_data = 12'b001110100111;
		16'b1011111000001110: color_data = 12'b001110100111;
		16'b1011111000001111: color_data = 12'b001110100111;
		16'b1011111000010000: color_data = 12'b001110100111;
		16'b1011111000010001: color_data = 12'b001110100111;
		16'b1011111000010010: color_data = 12'b001110100111;
		16'b1011111000010011: color_data = 12'b001110100111;
		16'b1011111000010100: color_data = 12'b001110100111;
		16'b1011111000010101: color_data = 12'b001110100111;
		16'b1011111000010110: color_data = 12'b001110100111;
		16'b1011111000010111: color_data = 12'b001110100111;
		16'b1011111000011000: color_data = 12'b001110100111;
		16'b1011111000011001: color_data = 12'b001110100111;
		16'b1011111000011010: color_data = 12'b001110100111;
		16'b1011111000011011: color_data = 12'b001110100111;
		16'b1011111000011100: color_data = 12'b001110100111;
		16'b1011111000011101: color_data = 12'b001110100111;
		16'b1011111000011110: color_data = 12'b001110100111;
		16'b1011111000011111: color_data = 12'b001110100111;
		16'b1011111000100000: color_data = 12'b001110100111;
		16'b1011111000100001: color_data = 12'b001110100111;
		16'b1011111000100010: color_data = 12'b001110100111;
		16'b1011111000100011: color_data = 12'b001110100111;
		16'b1011111000100100: color_data = 12'b001110100111;
		16'b1011111000101011: color_data = 12'b001110100111;
		16'b1011111000101100: color_data = 12'b001110100111;
		16'b1011111000101101: color_data = 12'b001110100111;
		16'b1011111000101110: color_data = 12'b001110100111;
		16'b1011111000101111: color_data = 12'b001110100111;
		16'b1011111000110000: color_data = 12'b001110100111;
		16'b1011111000110001: color_data = 12'b001110100111;
		16'b1011111000110010: color_data = 12'b001110100111;
		16'b1011111000110011: color_data = 12'b001110100111;
		16'b1011111000110100: color_data = 12'b001110100111;
		16'b1011111000110101: color_data = 12'b001110100111;
		16'b1011111000110110: color_data = 12'b001110100111;
		16'b1011111000110111: color_data = 12'b001110100111;
		16'b1011111001000100: color_data = 12'b001110100111;
		16'b1011111001000101: color_data = 12'b001110100111;
		16'b1011111001000110: color_data = 12'b001110100111;
		16'b1011111001000111: color_data = 12'b001110100111;
		16'b1011111001001000: color_data = 12'b001110100111;
		16'b1011111001001001: color_data = 12'b001110100111;
		16'b1011111001001010: color_data = 12'b001110100111;
		16'b1011111001001011: color_data = 12'b001110100111;
		16'b1011111001001100: color_data = 12'b001110100111;
		16'b1011111001001101: color_data = 12'b001110100111;
		16'b1011111001001110: color_data = 12'b001110100111;
		16'b1011111001001111: color_data = 12'b001110100111;
		16'b1011111001010110: color_data = 12'b001110100111;
		16'b1011111001010111: color_data = 12'b001110100111;
		16'b1011111001011000: color_data = 12'b001110100111;
		16'b1011111001011001: color_data = 12'b001110100111;
		16'b1011111001011010: color_data = 12'b001110100111;
		16'b1011111001011011: color_data = 12'b001110100111;
		16'b1011111001011100: color_data = 12'b001110100111;
		16'b1011111001011101: color_data = 12'b001110100111;
		16'b1011111001011110: color_data = 12'b001110100111;
		16'b1011111001011111: color_data = 12'b001110100111;
		16'b1011111001100000: color_data = 12'b001110100111;
		16'b1011111001100001: color_data = 12'b001110100111;
		16'b1011111001100010: color_data = 12'b001110100111;
		16'b1011111001100011: color_data = 12'b001110100111;
		16'b1011111001100100: color_data = 12'b001110100111;
		16'b1011111001100101: color_data = 12'b001110100111;
		16'b1011111001100110: color_data = 12'b001110100111;
		16'b1011111001100111: color_data = 12'b001110100111;
		16'b1011111001101000: color_data = 12'b001110100111;
		16'b1011111001101001: color_data = 12'b001110100111;
		16'b1011111001101010: color_data = 12'b001110100111;
		16'b1011111001101011: color_data = 12'b001110100111;
		16'b1011111001101100: color_data = 12'b001110100111;
		16'b1011111001101101: color_data = 12'b001110100111;
		16'b1011111001101110: color_data = 12'b001110100111;
		16'b1011111001110101: color_data = 12'b001110100111;
		16'b1011111001110110: color_data = 12'b001110100111;
		16'b1011111001110111: color_data = 12'b001110100111;
		16'b1011111001111000: color_data = 12'b001110100111;
		16'b1011111001111001: color_data = 12'b001110100111;
		16'b1011111001111010: color_data = 12'b001110100111;
		16'b1011111001111011: color_data = 12'b001110100111;
		16'b1011111001111100: color_data = 12'b001110100111;
		16'b1011111001111101: color_data = 12'b001110100111;
		16'b1011111001111110: color_data = 12'b001110100111;
		16'b1011111001111111: color_data = 12'b001110100111;
		16'b1011111010000000: color_data = 12'b001110100111;
		16'b1011111010001101: color_data = 12'b001110100111;
		16'b1011111010001110: color_data = 12'b001110100111;
		16'b1011111010001111: color_data = 12'b001110100111;
		16'b1011111010010000: color_data = 12'b001110100111;
		16'b1011111010010001: color_data = 12'b001110100111;
		16'b1011111010010010: color_data = 12'b001110100111;
		16'b1011111010010011: color_data = 12'b001110100111;
		16'b1011111010010100: color_data = 12'b001110100111;
		16'b1011111010010101: color_data = 12'b001110100111;
		16'b1011111010010110: color_data = 12'b001110100111;
		16'b1011111010010111: color_data = 12'b001110100111;
		16'b1011111010011000: color_data = 12'b001110100111;
		16'b1011111010011001: color_data = 12'b001110100111;
		16'b1011111010100000: color_data = 12'b001110100111;
		16'b1011111010100001: color_data = 12'b001110100111;
		16'b1011111010100010: color_data = 12'b001110100111;
		16'b1011111010100011: color_data = 12'b001110100111;
		16'b1011111010100100: color_data = 12'b001110100111;
		16'b1011111010100101: color_data = 12'b001110100111;
		16'b1011111010100110: color_data = 12'b001110100111;
		16'b1011111010100111: color_data = 12'b001110100111;
		16'b1011111010101000: color_data = 12'b001110100111;
		16'b1011111010101001: color_data = 12'b001110100111;
		16'b1011111010101010: color_data = 12'b001110100111;
		16'b1011111010101011: color_data = 12'b001110100111;
		16'b1011111010101100: color_data = 12'b001110100111;
		16'b1011111010101101: color_data = 12'b001110100111;
		16'b1011111010101110: color_data = 12'b001110100111;
		16'b1011111010101111: color_data = 12'b001110100111;
		16'b1011111010110000: color_data = 12'b001110100111;
		16'b1011111010110001: color_data = 12'b001110100111;
		16'b1011111010110010: color_data = 12'b001110100111;
		16'b1011111010110011: color_data = 12'b001110100111;
		16'b1011111010110100: color_data = 12'b001110100111;
		16'b1011111010110101: color_data = 12'b001110100111;
		16'b1011111010110110: color_data = 12'b001110100111;
		16'b1011111010110111: color_data = 12'b001110100111;
		16'b1011111010111000: color_data = 12'b001110100111;
		16'b1011111010111001: color_data = 12'b001110100111;
		16'b1011111010111010: color_data = 12'b001110100111;
		16'b1011111010111011: color_data = 12'b001110100111;
		16'b1011111010111100: color_data = 12'b001110100111;
		16'b1011111010111101: color_data = 12'b001110100111;
		16'b1011111010111110: color_data = 12'b001110100111;
		16'b1011111010111111: color_data = 12'b001110100111;
		16'b1011111011000000: color_data = 12'b001110100111;
		16'b1011111011000001: color_data = 12'b001110100111;
		16'b1011111011000010: color_data = 12'b001110100111;
		16'b1011111011000011: color_data = 12'b001110100111;
		16'b1011111011000100: color_data = 12'b001110100111;
		16'b1011111011001011: color_data = 12'b001110100111;
		16'b1011111011001100: color_data = 12'b001110100111;
		16'b1011111011001101: color_data = 12'b001110100111;
		16'b1011111011001110: color_data = 12'b001110100111;
		16'b1011111011001111: color_data = 12'b001110100111;
		16'b1011111011010000: color_data = 12'b001110100111;
		16'b1011111011010001: color_data = 12'b001110100111;
		16'b1011111011010010: color_data = 12'b001110100111;
		16'b1011111011010011: color_data = 12'b001110100111;
		16'b1011111011010100: color_data = 12'b001110100111;
		16'b1011111011010101: color_data = 12'b001110100111;
		16'b1011111011010110: color_data = 12'b001110100111;
		16'b1011111011111100: color_data = 12'b001110100111;
		16'b1011111011111101: color_data = 12'b001110100111;
		16'b1011111011111110: color_data = 12'b001110100111;
		16'b1011111011111111: color_data = 12'b001110100111;
		16'b1011111100000000: color_data = 12'b001110100111;
		16'b1011111100000001: color_data = 12'b001110100111;
		16'b1011111100000010: color_data = 12'b001110100111;
		16'b1011111100000011: color_data = 12'b001110100111;
		16'b1011111100000100: color_data = 12'b001110100111;
		16'b1011111100000101: color_data = 12'b001110100111;
		16'b1011111100000110: color_data = 12'b001110100111;
		16'b1011111100000111: color_data = 12'b001110100111;
		16'b1011111100001000: color_data = 12'b001110100111;
		16'b1011111100001001: color_data = 12'b001110100111;
		16'b1011111100001010: color_data = 12'b001110100111;
		16'b1011111100001011: color_data = 12'b001110100111;
		16'b1011111100001100: color_data = 12'b001110100111;
		16'b1011111100001101: color_data = 12'b001110100111;
		16'b1011111100001110: color_data = 12'b001110100111;
		16'b1011111100001111: color_data = 12'b001110100111;
		16'b1011111100010000: color_data = 12'b001110100111;
		16'b1011111100010001: color_data = 12'b001110100111;
		16'b1011111100010010: color_data = 12'b001110100111;
		16'b1011111100010011: color_data = 12'b001110100111;
		16'b1011111100010100: color_data = 12'b001110100111;
		16'b1011111100010101: color_data = 12'b001110100111;
		16'b1011111100010110: color_data = 12'b001110100111;
		16'b1011111100010111: color_data = 12'b001110100111;
		16'b1011111100011000: color_data = 12'b001110100111;
		16'b1011111100011001: color_data = 12'b001110100111;
		16'b1011111100011010: color_data = 12'b001110100111;
		16'b1011111100011011: color_data = 12'b001110100111;
		16'b1011111100011100: color_data = 12'b001110100111;
		16'b1011111100011101: color_data = 12'b001110100111;
		16'b1011111100011110: color_data = 12'b001110100111;
		16'b1011111100011111: color_data = 12'b001110100111;
		16'b1011111100100000: color_data = 12'b001110100111;
		16'b1011111100101101: color_data = 12'b001110100111;
		16'b1011111100101110: color_data = 12'b001110100111;
		16'b1011111100101111: color_data = 12'b001110100111;
		16'b1011111100110000: color_data = 12'b001110100111;
		16'b1011111100110001: color_data = 12'b001110100111;
		16'b1011111100110010: color_data = 12'b001110100111;
		16'b1011111100110011: color_data = 12'b001110100111;
		16'b1011111100110100: color_data = 12'b001110100111;
		16'b1011111100110101: color_data = 12'b001110100111;
		16'b1011111100110110: color_data = 12'b001110100111;
		16'b1011111100110111: color_data = 12'b001110100111;
		16'b1011111100111000: color_data = 12'b001110100111;
		16'b1011111101000101: color_data = 12'b001110100111;
		16'b1011111101000110: color_data = 12'b001110100111;
		16'b1011111101000111: color_data = 12'b001110100111;
		16'b1011111101001000: color_data = 12'b001110100111;
		16'b1011111101001001: color_data = 12'b001110100111;
		16'b1011111101001010: color_data = 12'b001110100111;
		16'b1011111101001011: color_data = 12'b001110100111;
		16'b1011111101001100: color_data = 12'b001110100111;
		16'b1011111101001101: color_data = 12'b001110100111;
		16'b1011111101001110: color_data = 12'b001110100111;
		16'b1011111101001111: color_data = 12'b001110100111;
		16'b1011111101010000: color_data = 12'b001110100111;
		16'b1011111101010001: color_data = 12'b001110100111;
		16'b1011111101011000: color_data = 12'b001110100111;
		16'b1011111101011001: color_data = 12'b001110100111;
		16'b1011111101011010: color_data = 12'b001110100111;
		16'b1011111101011011: color_data = 12'b001110100111;
		16'b1011111101011100: color_data = 12'b001110100111;
		16'b1011111101011101: color_data = 12'b001110100111;
		16'b1011111101011110: color_data = 12'b001110100111;
		16'b1011111101011111: color_data = 12'b001110100111;
		16'b1011111101100000: color_data = 12'b001110100111;
		16'b1011111101100001: color_data = 12'b001110100111;
		16'b1011111101100010: color_data = 12'b001110100111;
		16'b1011111101100011: color_data = 12'b001110100111;
		16'b1011111101100100: color_data = 12'b001110100111;
		16'b1011111101100101: color_data = 12'b001110100111;
		16'b1011111101100110: color_data = 12'b001110100111;
		16'b1011111101100111: color_data = 12'b001110100111;
		16'b1011111101101000: color_data = 12'b001110100111;
		16'b1011111101101001: color_data = 12'b001110100111;
		16'b1011111101101010: color_data = 12'b001110100111;
		16'b1011111101101011: color_data = 12'b001110100111;
		16'b1011111101101100: color_data = 12'b001110100111;
		16'b1011111101101101: color_data = 12'b001110100111;
		16'b1011111101101110: color_data = 12'b001110100111;
		16'b1011111101101111: color_data = 12'b001110100111;
		16'b1011111101110000: color_data = 12'b001110100111;
		16'b1011111101110001: color_data = 12'b001110100111;
		16'b1011111101110010: color_data = 12'b001110100111;
		16'b1011111101110011: color_data = 12'b001110100111;
		16'b1011111101110100: color_data = 12'b001110100111;
		16'b1011111101110101: color_data = 12'b001110100111;
		16'b1011111101110110: color_data = 12'b001110100111;
		16'b1011111101110111: color_data = 12'b001110100111;
		16'b1011111101111000: color_data = 12'b001110100111;
		16'b1011111101111001: color_data = 12'b001110100111;
		16'b1011111101111010: color_data = 12'b001110100111;
		16'b1011111101111011: color_data = 12'b001110100111;
		16'b1100000000000000: color_data = 12'b001110100111;
		16'b1100000000000001: color_data = 12'b001110100111;
		16'b1100000000000010: color_data = 12'b001110100111;
		16'b1100000000000011: color_data = 12'b001110100111;
		16'b1100000000000100: color_data = 12'b001110100111;
		16'b1100000000000101: color_data = 12'b001110100111;
		16'b1100000000000110: color_data = 12'b001110100111;
		16'b1100000000000111: color_data = 12'b001110100111;
		16'b1100000000001000: color_data = 12'b001110100111;
		16'b1100000000001001: color_data = 12'b001110100111;
		16'b1100000000001010: color_data = 12'b001110100111;
		16'b1100000000001011: color_data = 12'b001110100111;
		16'b1100000000001100: color_data = 12'b001110100111;
		16'b1100000000001101: color_data = 12'b001110100111;
		16'b1100000000001110: color_data = 12'b001110100111;
		16'b1100000000001111: color_data = 12'b001110100111;
		16'b1100000000010000: color_data = 12'b001110100111;
		16'b1100000000010001: color_data = 12'b001110100111;
		16'b1100000000010010: color_data = 12'b001110100111;
		16'b1100000000010011: color_data = 12'b001110100111;
		16'b1100000000010100: color_data = 12'b001110100111;
		16'b1100000000010101: color_data = 12'b001110100111;
		16'b1100000000010110: color_data = 12'b001110100111;
		16'b1100000000010111: color_data = 12'b001110100111;
		16'b1100000000011000: color_data = 12'b001110100111;
		16'b1100000000011001: color_data = 12'b001110100111;
		16'b1100000000011010: color_data = 12'b001110100111;
		16'b1100000000011011: color_data = 12'b001110100111;
		16'b1100000000011100: color_data = 12'b001110100111;
		16'b1100000000011101: color_data = 12'b001110100111;
		16'b1100000000011110: color_data = 12'b001110100111;
		16'b1100000000011111: color_data = 12'b001110100111;
		16'b1100000000100000: color_data = 12'b001110100111;
		16'b1100000000100001: color_data = 12'b001110100111;
		16'b1100000000100010: color_data = 12'b001110100111;
		16'b1100000000100011: color_data = 12'b001110100111;
		16'b1100000000100100: color_data = 12'b001110100111;
		16'b1100000000101011: color_data = 12'b001110100111;
		16'b1100000000101100: color_data = 12'b001110100111;
		16'b1100000000101101: color_data = 12'b001110100111;
		16'b1100000000101110: color_data = 12'b001110100111;
		16'b1100000000101111: color_data = 12'b001110100111;
		16'b1100000000110000: color_data = 12'b001110100111;
		16'b1100000000110001: color_data = 12'b001110100111;
		16'b1100000000110010: color_data = 12'b001110100111;
		16'b1100000000110011: color_data = 12'b001110100111;
		16'b1100000000110100: color_data = 12'b001110100111;
		16'b1100000000110101: color_data = 12'b001110100111;
		16'b1100000000110110: color_data = 12'b001110100111;
		16'b1100000000110111: color_data = 12'b001110100111;
		16'b1100000001000100: color_data = 12'b001110100111;
		16'b1100000001000101: color_data = 12'b001110100111;
		16'b1100000001000110: color_data = 12'b001110100111;
		16'b1100000001000111: color_data = 12'b001110100111;
		16'b1100000001001000: color_data = 12'b001110100111;
		16'b1100000001001001: color_data = 12'b001110100111;
		16'b1100000001001010: color_data = 12'b001110100111;
		16'b1100000001001011: color_data = 12'b001110100111;
		16'b1100000001001100: color_data = 12'b001110100111;
		16'b1100000001001101: color_data = 12'b001110100111;
		16'b1100000001001110: color_data = 12'b001110100111;
		16'b1100000001001111: color_data = 12'b001110100111;
		16'b1100000001010110: color_data = 12'b001110100111;
		16'b1100000001010111: color_data = 12'b001110100111;
		16'b1100000001011000: color_data = 12'b001110100111;
		16'b1100000001011001: color_data = 12'b001110100111;
		16'b1100000001011010: color_data = 12'b001110100111;
		16'b1100000001011011: color_data = 12'b001110100111;
		16'b1100000001011100: color_data = 12'b001110100111;
		16'b1100000001011101: color_data = 12'b001110100111;
		16'b1100000001011110: color_data = 12'b001110100111;
		16'b1100000001011111: color_data = 12'b001110100111;
		16'b1100000001100000: color_data = 12'b001110100111;
		16'b1100000001100001: color_data = 12'b001110100111;
		16'b1100000001100010: color_data = 12'b001110100111;
		16'b1100000001100011: color_data = 12'b001110100111;
		16'b1100000001100100: color_data = 12'b001110100111;
		16'b1100000001100101: color_data = 12'b001110100111;
		16'b1100000001100110: color_data = 12'b001110100111;
		16'b1100000001100111: color_data = 12'b001110100111;
		16'b1100000001101000: color_data = 12'b001110100111;
		16'b1100000001101001: color_data = 12'b001110100111;
		16'b1100000001101010: color_data = 12'b001110100111;
		16'b1100000001101011: color_data = 12'b001110100111;
		16'b1100000001101100: color_data = 12'b001110100111;
		16'b1100000001101101: color_data = 12'b001110100111;
		16'b1100000001101110: color_data = 12'b001110100111;
		16'b1100000001110101: color_data = 12'b001110100111;
		16'b1100000001110110: color_data = 12'b001110100111;
		16'b1100000001110111: color_data = 12'b001110100111;
		16'b1100000001111000: color_data = 12'b001110100111;
		16'b1100000001111001: color_data = 12'b001110100111;
		16'b1100000001111010: color_data = 12'b001110100111;
		16'b1100000001111011: color_data = 12'b001110100111;
		16'b1100000001111100: color_data = 12'b001110100111;
		16'b1100000001111101: color_data = 12'b001110100111;
		16'b1100000001111110: color_data = 12'b001110100111;
		16'b1100000001111111: color_data = 12'b001110100111;
		16'b1100000010000000: color_data = 12'b001110100111;
		16'b1100000010001101: color_data = 12'b001110100111;
		16'b1100000010001110: color_data = 12'b001110100111;
		16'b1100000010001111: color_data = 12'b001110100111;
		16'b1100000010010000: color_data = 12'b001110100111;
		16'b1100000010010001: color_data = 12'b001110100111;
		16'b1100000010010010: color_data = 12'b001110100111;
		16'b1100000010010011: color_data = 12'b001110100111;
		16'b1100000010010100: color_data = 12'b001110100111;
		16'b1100000010010101: color_data = 12'b001110100111;
		16'b1100000010010110: color_data = 12'b001110100111;
		16'b1100000010010111: color_data = 12'b001110100111;
		16'b1100000010011000: color_data = 12'b001110100111;
		16'b1100000010011001: color_data = 12'b001110100111;
		16'b1100000010100000: color_data = 12'b001110100111;
		16'b1100000010100001: color_data = 12'b001110100111;
		16'b1100000010100010: color_data = 12'b001110100111;
		16'b1100000010100011: color_data = 12'b001110100111;
		16'b1100000010100100: color_data = 12'b001110100111;
		16'b1100000010100101: color_data = 12'b001110100111;
		16'b1100000010100110: color_data = 12'b001110100111;
		16'b1100000010100111: color_data = 12'b001110100111;
		16'b1100000010101000: color_data = 12'b001110100111;
		16'b1100000010101001: color_data = 12'b001110100111;
		16'b1100000010101010: color_data = 12'b001110100111;
		16'b1100000010101011: color_data = 12'b001110100111;
		16'b1100000010101100: color_data = 12'b001110100111;
		16'b1100000010101101: color_data = 12'b001110100111;
		16'b1100000010101110: color_data = 12'b001110100111;
		16'b1100000010101111: color_data = 12'b001110100111;
		16'b1100000010110000: color_data = 12'b001110100111;
		16'b1100000010110001: color_data = 12'b001110100111;
		16'b1100000010110010: color_data = 12'b001110100111;
		16'b1100000010110011: color_data = 12'b001110100111;
		16'b1100000010110100: color_data = 12'b001110100111;
		16'b1100000010110101: color_data = 12'b001110100111;
		16'b1100000010110110: color_data = 12'b001110100111;
		16'b1100000010110111: color_data = 12'b001110100111;
		16'b1100000010111000: color_data = 12'b001110100111;
		16'b1100000010111001: color_data = 12'b001110100111;
		16'b1100000010111010: color_data = 12'b001110100111;
		16'b1100000010111011: color_data = 12'b001110100111;
		16'b1100000010111100: color_data = 12'b001110100111;
		16'b1100000010111101: color_data = 12'b001110100111;
		16'b1100000010111110: color_data = 12'b001110100111;
		16'b1100000010111111: color_data = 12'b001110100111;
		16'b1100000011000000: color_data = 12'b001110100111;
		16'b1100000011000001: color_data = 12'b001110100111;
		16'b1100000011000010: color_data = 12'b001110100111;
		16'b1100000011000011: color_data = 12'b001110100111;
		16'b1100000011000100: color_data = 12'b001110100111;
		16'b1100000011001011: color_data = 12'b001110100111;
		16'b1100000011001100: color_data = 12'b001110100111;
		16'b1100000011001101: color_data = 12'b001110100111;
		16'b1100000011001110: color_data = 12'b001110100111;
		16'b1100000011001111: color_data = 12'b001110100111;
		16'b1100000011010000: color_data = 12'b001110100111;
		16'b1100000011010001: color_data = 12'b001110100111;
		16'b1100000011010010: color_data = 12'b001110100111;
		16'b1100000011010011: color_data = 12'b001110100111;
		16'b1100000011010100: color_data = 12'b001110100111;
		16'b1100000011010101: color_data = 12'b001110100111;
		16'b1100000011010110: color_data = 12'b001110100111;
		16'b1100000011111100: color_data = 12'b001110100111;
		16'b1100000011111101: color_data = 12'b001110100111;
		16'b1100000011111110: color_data = 12'b001110100111;
		16'b1100000011111111: color_data = 12'b001110100111;
		16'b1100000100000000: color_data = 12'b001110100111;
		16'b1100000100000001: color_data = 12'b001110100111;
		16'b1100000100000010: color_data = 12'b001110100111;
		16'b1100000100000011: color_data = 12'b001110100111;
		16'b1100000100000100: color_data = 12'b001110100111;
		16'b1100000100000101: color_data = 12'b001110100111;
		16'b1100000100000110: color_data = 12'b001110100111;
		16'b1100000100000111: color_data = 12'b001110100111;
		16'b1100000100001000: color_data = 12'b001110100111;
		16'b1100000100001001: color_data = 12'b001110100111;
		16'b1100000100001010: color_data = 12'b001110100111;
		16'b1100000100001011: color_data = 12'b001110100111;
		16'b1100000100001100: color_data = 12'b001110100111;
		16'b1100000100001101: color_data = 12'b001110100111;
		16'b1100000100001110: color_data = 12'b001110100111;
		16'b1100000100001111: color_data = 12'b001110100111;
		16'b1100000100010000: color_data = 12'b001110100111;
		16'b1100000100010001: color_data = 12'b001110100111;
		16'b1100000100010010: color_data = 12'b001110100111;
		16'b1100000100010011: color_data = 12'b001110100111;
		16'b1100000100010100: color_data = 12'b001110100111;
		16'b1100000100010101: color_data = 12'b001110100111;
		16'b1100000100010110: color_data = 12'b001110100111;
		16'b1100000100010111: color_data = 12'b001110100111;
		16'b1100000100011000: color_data = 12'b001110100111;
		16'b1100000100011001: color_data = 12'b001110100111;
		16'b1100000100011010: color_data = 12'b001110100111;
		16'b1100000100011011: color_data = 12'b001110100111;
		16'b1100000100011100: color_data = 12'b001110100111;
		16'b1100000100011101: color_data = 12'b001110100111;
		16'b1100000100011110: color_data = 12'b001110100111;
		16'b1100000100011111: color_data = 12'b001110100111;
		16'b1100000100100000: color_data = 12'b001110100111;
		16'b1100000100101101: color_data = 12'b001110100111;
		16'b1100000100101110: color_data = 12'b001110100111;
		16'b1100000100101111: color_data = 12'b001110100111;
		16'b1100000100110000: color_data = 12'b001110100111;
		16'b1100000100110001: color_data = 12'b001110100111;
		16'b1100000100110010: color_data = 12'b001110100111;
		16'b1100000100110011: color_data = 12'b001110100111;
		16'b1100000100110100: color_data = 12'b001110100111;
		16'b1100000100110101: color_data = 12'b001110100111;
		16'b1100000100110110: color_data = 12'b001110100111;
		16'b1100000100110111: color_data = 12'b001110100111;
		16'b1100000100111000: color_data = 12'b001110100111;
		16'b1100000101000101: color_data = 12'b001110100111;
		16'b1100000101000110: color_data = 12'b001110100111;
		16'b1100000101000111: color_data = 12'b001110100111;
		16'b1100000101001000: color_data = 12'b001110100111;
		16'b1100000101001001: color_data = 12'b001110100111;
		16'b1100000101001010: color_data = 12'b001110100111;
		16'b1100000101001011: color_data = 12'b001110100111;
		16'b1100000101001100: color_data = 12'b001110100111;
		16'b1100000101001101: color_data = 12'b001110100111;
		16'b1100000101001110: color_data = 12'b001110100111;
		16'b1100000101001111: color_data = 12'b001110100111;
		16'b1100000101010000: color_data = 12'b001110100111;
		16'b1100000101010001: color_data = 12'b001110100111;
		16'b1100000101011000: color_data = 12'b001110100111;
		16'b1100000101011001: color_data = 12'b001110100111;
		16'b1100000101011010: color_data = 12'b001110100111;
		16'b1100000101011011: color_data = 12'b001110100111;
		16'b1100000101011100: color_data = 12'b001110100111;
		16'b1100000101011101: color_data = 12'b001110100111;
		16'b1100000101011110: color_data = 12'b001110100111;
		16'b1100000101011111: color_data = 12'b001110100111;
		16'b1100000101100000: color_data = 12'b001110100111;
		16'b1100000101100001: color_data = 12'b001110100111;
		16'b1100000101100010: color_data = 12'b001110100111;
		16'b1100000101100011: color_data = 12'b001110100111;
		16'b1100000101100100: color_data = 12'b001110100111;
		16'b1100000101100101: color_data = 12'b001110100111;
		16'b1100000101100110: color_data = 12'b001110100111;
		16'b1100000101100111: color_data = 12'b001110100111;
		16'b1100000101101000: color_data = 12'b001110100111;
		16'b1100000101101001: color_data = 12'b001110100111;
		16'b1100000101101010: color_data = 12'b001110100111;
		16'b1100000101101011: color_data = 12'b001110100111;
		16'b1100000101101100: color_data = 12'b001110100111;
		16'b1100000101101101: color_data = 12'b001110100111;
		16'b1100000101101110: color_data = 12'b001110100111;
		16'b1100000101101111: color_data = 12'b001110100111;
		16'b1100000101110000: color_data = 12'b001110100111;
		16'b1100000101110001: color_data = 12'b001110100111;
		16'b1100000101110010: color_data = 12'b001110100111;
		16'b1100000101110011: color_data = 12'b001110100111;
		16'b1100000101110100: color_data = 12'b001110100111;
		16'b1100000101110101: color_data = 12'b001110100111;
		16'b1100000101110110: color_data = 12'b001110100111;
		16'b1100000101110111: color_data = 12'b001110100111;
		16'b1100000101111000: color_data = 12'b001110100111;
		16'b1100000101111001: color_data = 12'b001110100111;
		16'b1100000101111010: color_data = 12'b001110100111;
		16'b1100000101111011: color_data = 12'b001110100111;
		16'b1100001000000000: color_data = 12'b001110100111;
		16'b1100001000000001: color_data = 12'b001110100111;
		16'b1100001000000010: color_data = 12'b001110100111;
		16'b1100001000000011: color_data = 12'b001110100111;
		16'b1100001000000100: color_data = 12'b001110100111;
		16'b1100001000000101: color_data = 12'b001110100111;
		16'b1100001000000110: color_data = 12'b001110100111;
		16'b1100001000000111: color_data = 12'b001110100111;
		16'b1100001000001000: color_data = 12'b001110100111;
		16'b1100001000001001: color_data = 12'b001110100111;
		16'b1100001000001010: color_data = 12'b001110100111;
		16'b1100001000001011: color_data = 12'b001110100111;
		16'b1100001000001100: color_data = 12'b001110100111;
		16'b1100001000001101: color_data = 12'b001110100111;
		16'b1100001000001110: color_data = 12'b001110100111;
		16'b1100001000001111: color_data = 12'b001110100111;
		16'b1100001000010000: color_data = 12'b001110100111;
		16'b1100001000010001: color_data = 12'b001110100111;
		16'b1100001000010010: color_data = 12'b001110100111;
		16'b1100001000010011: color_data = 12'b001110100111;
		16'b1100001000010100: color_data = 12'b001110100111;
		16'b1100001000010101: color_data = 12'b001110100111;
		16'b1100001000010110: color_data = 12'b001110100111;
		16'b1100001000010111: color_data = 12'b001110100111;
		16'b1100001000011000: color_data = 12'b001110100111;
		16'b1100001000011001: color_data = 12'b001110100111;
		16'b1100001000011010: color_data = 12'b001110100111;
		16'b1100001000011011: color_data = 12'b001110100111;
		16'b1100001000011100: color_data = 12'b001110100111;
		16'b1100001000011101: color_data = 12'b001110100111;
		16'b1100001000011110: color_data = 12'b001110100111;
		16'b1100001000011111: color_data = 12'b001110100111;
		16'b1100001000100000: color_data = 12'b001110100111;
		16'b1100001000100001: color_data = 12'b001110100111;
		16'b1100001000100010: color_data = 12'b001110100111;
		16'b1100001000100011: color_data = 12'b001110100111;
		16'b1100001000100100: color_data = 12'b001110100111;
		16'b1100001000101011: color_data = 12'b001110100111;
		16'b1100001000101100: color_data = 12'b001110100111;
		16'b1100001000101101: color_data = 12'b001110100111;
		16'b1100001000101110: color_data = 12'b001110100111;
		16'b1100001000101111: color_data = 12'b001110100111;
		16'b1100001000110000: color_data = 12'b001110100111;
		16'b1100001000110001: color_data = 12'b001110100111;
		16'b1100001000110010: color_data = 12'b001110100111;
		16'b1100001000110011: color_data = 12'b001110100111;
		16'b1100001000110100: color_data = 12'b001110100111;
		16'b1100001000110101: color_data = 12'b001110100111;
		16'b1100001000110110: color_data = 12'b001110100111;
		16'b1100001000110111: color_data = 12'b001110100111;
		16'b1100001001000100: color_data = 12'b001110100111;
		16'b1100001001000101: color_data = 12'b001110100111;
		16'b1100001001000110: color_data = 12'b001110100111;
		16'b1100001001000111: color_data = 12'b001110100111;
		16'b1100001001001000: color_data = 12'b001110100111;
		16'b1100001001001001: color_data = 12'b001110100111;
		16'b1100001001001010: color_data = 12'b001110100111;
		16'b1100001001001011: color_data = 12'b001110100111;
		16'b1100001001001100: color_data = 12'b001110100111;
		16'b1100001001001101: color_data = 12'b001110100111;
		16'b1100001001001110: color_data = 12'b001110100111;
		16'b1100001001001111: color_data = 12'b001110100111;
		16'b1100001001010110: color_data = 12'b001110100111;
		16'b1100001001010111: color_data = 12'b001110100111;
		16'b1100001001011000: color_data = 12'b001110100111;
		16'b1100001001011001: color_data = 12'b001110100111;
		16'b1100001001011010: color_data = 12'b001110100111;
		16'b1100001001011011: color_data = 12'b001110100111;
		16'b1100001001011100: color_data = 12'b001110100111;
		16'b1100001001011101: color_data = 12'b001110100111;
		16'b1100001001011110: color_data = 12'b001110100111;
		16'b1100001001011111: color_data = 12'b001110100111;
		16'b1100001001100000: color_data = 12'b001110100111;
		16'b1100001001100001: color_data = 12'b001110100111;
		16'b1100001001100010: color_data = 12'b001110100111;
		16'b1100001001100011: color_data = 12'b001110100111;
		16'b1100001001100100: color_data = 12'b001110100111;
		16'b1100001001100101: color_data = 12'b001110100111;
		16'b1100001001100110: color_data = 12'b001110100111;
		16'b1100001001100111: color_data = 12'b001110100111;
		16'b1100001001101000: color_data = 12'b001110100111;
		16'b1100001001101001: color_data = 12'b001110100111;
		16'b1100001001101010: color_data = 12'b001110100111;
		16'b1100001001101011: color_data = 12'b001110100111;
		16'b1100001001101100: color_data = 12'b001110100111;
		16'b1100001001101101: color_data = 12'b001110100111;
		16'b1100001001101110: color_data = 12'b001110100111;
		16'b1100001001110101: color_data = 12'b001110100111;
		16'b1100001001110110: color_data = 12'b001110100111;
		16'b1100001001110111: color_data = 12'b001110100111;
		16'b1100001001111000: color_data = 12'b001110100111;
		16'b1100001001111001: color_data = 12'b001110100111;
		16'b1100001001111010: color_data = 12'b001110100111;
		16'b1100001001111011: color_data = 12'b001110100111;
		16'b1100001001111100: color_data = 12'b001110100111;
		16'b1100001001111101: color_data = 12'b001110100111;
		16'b1100001001111110: color_data = 12'b001110100111;
		16'b1100001001111111: color_data = 12'b001110100111;
		16'b1100001010000000: color_data = 12'b001110100111;
		16'b1100001010001101: color_data = 12'b001110100111;
		16'b1100001010001110: color_data = 12'b001110100111;
		16'b1100001010001111: color_data = 12'b001110100111;
		16'b1100001010010000: color_data = 12'b001110100111;
		16'b1100001010010001: color_data = 12'b001110100111;
		16'b1100001010010010: color_data = 12'b001110100111;
		16'b1100001010010011: color_data = 12'b001110100111;
		16'b1100001010010100: color_data = 12'b001110100111;
		16'b1100001010010101: color_data = 12'b001110100111;
		16'b1100001010010110: color_data = 12'b001110100111;
		16'b1100001010010111: color_data = 12'b001110100111;
		16'b1100001010011000: color_data = 12'b001110100111;
		16'b1100001010011001: color_data = 12'b001110100111;
		16'b1100001010100000: color_data = 12'b001110100111;
		16'b1100001010100001: color_data = 12'b001110100111;
		16'b1100001010100010: color_data = 12'b001110100111;
		16'b1100001010100011: color_data = 12'b001110100111;
		16'b1100001010100100: color_data = 12'b001110100111;
		16'b1100001010100101: color_data = 12'b001110100111;
		16'b1100001010100110: color_data = 12'b001110100111;
		16'b1100001010100111: color_data = 12'b001110100111;
		16'b1100001010101000: color_data = 12'b001110100111;
		16'b1100001010101001: color_data = 12'b001110100111;
		16'b1100001010101010: color_data = 12'b001110100111;
		16'b1100001010101011: color_data = 12'b001110100111;
		16'b1100001010101100: color_data = 12'b001110100111;
		16'b1100001010101101: color_data = 12'b001110100111;
		16'b1100001010101110: color_data = 12'b001110100111;
		16'b1100001010101111: color_data = 12'b001110100111;
		16'b1100001010110000: color_data = 12'b001110100111;
		16'b1100001010110001: color_data = 12'b001110100111;
		16'b1100001010110010: color_data = 12'b001110100111;
		16'b1100001010110011: color_data = 12'b001110100111;
		16'b1100001010110100: color_data = 12'b001110100111;
		16'b1100001010110101: color_data = 12'b001110100111;
		16'b1100001010110110: color_data = 12'b001110100111;
		16'b1100001010110111: color_data = 12'b001110100111;
		16'b1100001010111000: color_data = 12'b001110100111;
		16'b1100001010111001: color_data = 12'b001110100111;
		16'b1100001010111010: color_data = 12'b001110100111;
		16'b1100001010111011: color_data = 12'b001110100111;
		16'b1100001010111100: color_data = 12'b001110100111;
		16'b1100001010111101: color_data = 12'b001110100111;
		16'b1100001010111110: color_data = 12'b001110100111;
		16'b1100001010111111: color_data = 12'b001110100111;
		16'b1100001011000000: color_data = 12'b001110100111;
		16'b1100001011000001: color_data = 12'b001110100111;
		16'b1100001011000010: color_data = 12'b001110100111;
		16'b1100001011000011: color_data = 12'b001110100111;
		16'b1100001011000100: color_data = 12'b001110100111;
		16'b1100001011001011: color_data = 12'b001110100111;
		16'b1100001011001100: color_data = 12'b001110100111;
		16'b1100001011001101: color_data = 12'b001110100111;
		16'b1100001011001110: color_data = 12'b001110100111;
		16'b1100001011001111: color_data = 12'b001110100111;
		16'b1100001011010000: color_data = 12'b001110100111;
		16'b1100001011010001: color_data = 12'b001110100111;
		16'b1100001011010010: color_data = 12'b001110100111;
		16'b1100001011010011: color_data = 12'b001110100111;
		16'b1100001011010100: color_data = 12'b001110100111;
		16'b1100001011010101: color_data = 12'b001110100111;
		16'b1100001011010110: color_data = 12'b001110100111;
		16'b1100001011111100: color_data = 12'b001110100111;
		16'b1100001011111101: color_data = 12'b001110100111;
		16'b1100001011111110: color_data = 12'b001110100111;
		16'b1100001011111111: color_data = 12'b001110100111;
		16'b1100001100000000: color_data = 12'b001110100111;
		16'b1100001100000001: color_data = 12'b001110100111;
		16'b1100001100000010: color_data = 12'b001110100111;
		16'b1100001100000011: color_data = 12'b001110100111;
		16'b1100001100000100: color_data = 12'b001110100111;
		16'b1100001100000101: color_data = 12'b001110100111;
		16'b1100001100000110: color_data = 12'b001110100111;
		16'b1100001100000111: color_data = 12'b001110100111;
		16'b1100001100001000: color_data = 12'b001110100111;
		16'b1100001100001001: color_data = 12'b001110100111;
		16'b1100001100001010: color_data = 12'b001110100111;
		16'b1100001100001011: color_data = 12'b001110100111;
		16'b1100001100001100: color_data = 12'b001110100111;
		16'b1100001100001101: color_data = 12'b001110100111;
		16'b1100001100001110: color_data = 12'b001110100111;
		16'b1100001100001111: color_data = 12'b001110100111;
		16'b1100001100010000: color_data = 12'b001110100111;
		16'b1100001100010001: color_data = 12'b001110100111;
		16'b1100001100010010: color_data = 12'b001110100111;
		16'b1100001100010011: color_data = 12'b001110100111;
		16'b1100001100010100: color_data = 12'b001110100111;
		16'b1100001100010101: color_data = 12'b001110100111;
		16'b1100001100010110: color_data = 12'b001110100111;
		16'b1100001100010111: color_data = 12'b001110100111;
		16'b1100001100011000: color_data = 12'b001110100111;
		16'b1100001100011001: color_data = 12'b001110100111;
		16'b1100001100011010: color_data = 12'b001110100111;
		16'b1100001100011011: color_data = 12'b001110100111;
		16'b1100001100011100: color_data = 12'b001110100111;
		16'b1100001100011101: color_data = 12'b001110100111;
		16'b1100001100011110: color_data = 12'b001110100111;
		16'b1100001100011111: color_data = 12'b001110100111;
		16'b1100001100100000: color_data = 12'b001110100111;
		16'b1100001100101101: color_data = 12'b001110100111;
		16'b1100001100101110: color_data = 12'b001110100111;
		16'b1100001100101111: color_data = 12'b001110100111;
		16'b1100001100110000: color_data = 12'b001110100111;
		16'b1100001100110001: color_data = 12'b001110100111;
		16'b1100001100110010: color_data = 12'b001110100111;
		16'b1100001100110011: color_data = 12'b001110100111;
		16'b1100001100110100: color_data = 12'b001110100111;
		16'b1100001100110101: color_data = 12'b001110100111;
		16'b1100001100110110: color_data = 12'b001110100111;
		16'b1100001100110111: color_data = 12'b001110100111;
		16'b1100001100111000: color_data = 12'b001110100111;
		16'b1100001101000101: color_data = 12'b001110100111;
		16'b1100001101000110: color_data = 12'b001110100111;
		16'b1100001101000111: color_data = 12'b001110100111;
		16'b1100001101001000: color_data = 12'b001110100111;
		16'b1100001101001001: color_data = 12'b001110100111;
		16'b1100001101001010: color_data = 12'b001110100111;
		16'b1100001101001011: color_data = 12'b001110100111;
		16'b1100001101001100: color_data = 12'b001110100111;
		16'b1100001101001101: color_data = 12'b001110100111;
		16'b1100001101001110: color_data = 12'b001110100111;
		16'b1100001101001111: color_data = 12'b001110100111;
		16'b1100001101010000: color_data = 12'b001110100111;
		16'b1100001101010001: color_data = 12'b001110100111;
		16'b1100001101011000: color_data = 12'b001110100111;
		16'b1100001101011001: color_data = 12'b001110100111;
		16'b1100001101011010: color_data = 12'b001110100111;
		16'b1100001101011011: color_data = 12'b001110100111;
		16'b1100001101011100: color_data = 12'b001110100111;
		16'b1100001101011101: color_data = 12'b001110100111;
		16'b1100001101011110: color_data = 12'b001110100111;
		16'b1100001101011111: color_data = 12'b001110100111;
		16'b1100001101100000: color_data = 12'b001110100111;
		16'b1100001101100001: color_data = 12'b001110100111;
		16'b1100001101100010: color_data = 12'b001110100111;
		16'b1100001101100011: color_data = 12'b001110100111;
		16'b1100001101100100: color_data = 12'b001110100111;
		16'b1100001101100101: color_data = 12'b001110100111;
		16'b1100001101100110: color_data = 12'b001110100111;
		16'b1100001101100111: color_data = 12'b001110100111;
		16'b1100001101101000: color_data = 12'b001110100111;
		16'b1100001101101001: color_data = 12'b001110100111;
		16'b1100001101101010: color_data = 12'b001110100111;
		16'b1100001101101011: color_data = 12'b001110100111;
		16'b1100001101101100: color_data = 12'b001110100111;
		16'b1100001101101101: color_data = 12'b001110100111;
		16'b1100001101101110: color_data = 12'b001110100111;
		16'b1100001101101111: color_data = 12'b001110100111;
		16'b1100001101110000: color_data = 12'b001110100111;
		16'b1100001101110001: color_data = 12'b001110100111;
		16'b1100001101110010: color_data = 12'b001110100111;
		16'b1100001101110011: color_data = 12'b001110100111;
		16'b1100001101110100: color_data = 12'b001110100111;
		16'b1100001101110101: color_data = 12'b001110100111;
		16'b1100001101110110: color_data = 12'b001110100111;
		16'b1100001101110111: color_data = 12'b001110100111;
		16'b1100001101111000: color_data = 12'b001110100111;
		16'b1100001101111001: color_data = 12'b001110100111;
		16'b1100001101111010: color_data = 12'b001110100111;
		16'b1100001101111011: color_data = 12'b001110100111;
		16'b1100010000000000: color_data = 12'b001110100111;
		16'b1100010000000001: color_data = 12'b001110100111;
		16'b1100010000000010: color_data = 12'b001110100111;
		16'b1100010000000011: color_data = 12'b001110100111;
		16'b1100010000000100: color_data = 12'b001110100111;
		16'b1100010000000101: color_data = 12'b001110100111;
		16'b1100010000000110: color_data = 12'b001110100111;
		16'b1100010000000111: color_data = 12'b001110100111;
		16'b1100010000001000: color_data = 12'b001110100111;
		16'b1100010000001001: color_data = 12'b001110100111;
		16'b1100010000001010: color_data = 12'b001110100111;
		16'b1100010000001011: color_data = 12'b001110100111;
		16'b1100010000001100: color_data = 12'b001110100111;
		16'b1100010000001101: color_data = 12'b001110100111;
		16'b1100010000001110: color_data = 12'b001110100111;
		16'b1100010000001111: color_data = 12'b001110100111;
		16'b1100010000010000: color_data = 12'b001110100111;
		16'b1100010000010001: color_data = 12'b001110100111;
		16'b1100010000010010: color_data = 12'b001110100111;
		16'b1100010000010011: color_data = 12'b001110100111;
		16'b1100010000010100: color_data = 12'b001110100111;
		16'b1100010000010101: color_data = 12'b001110100111;
		16'b1100010000010110: color_data = 12'b001110100111;
		16'b1100010000010111: color_data = 12'b001110100111;
		16'b1100010000011000: color_data = 12'b001110100111;
		16'b1100010000011001: color_data = 12'b001110100111;
		16'b1100010000011010: color_data = 12'b001110100111;
		16'b1100010000011011: color_data = 12'b001110100111;
		16'b1100010000011100: color_data = 12'b001110100111;
		16'b1100010000011101: color_data = 12'b001110100111;
		16'b1100010000011110: color_data = 12'b001110100111;
		16'b1100010000011111: color_data = 12'b001110100111;
		16'b1100010000100000: color_data = 12'b001110100111;
		16'b1100010000100001: color_data = 12'b001110100111;
		16'b1100010000100010: color_data = 12'b001110100111;
		16'b1100010000100011: color_data = 12'b001110100111;
		16'b1100010000100100: color_data = 12'b001110100111;
		16'b1100010000101011: color_data = 12'b001110100111;
		16'b1100010000101100: color_data = 12'b001110100111;
		16'b1100010000101101: color_data = 12'b001110100111;
		16'b1100010000101110: color_data = 12'b001110100111;
		16'b1100010000101111: color_data = 12'b001110100111;
		16'b1100010000110000: color_data = 12'b001110100111;
		16'b1100010000110001: color_data = 12'b001110100111;
		16'b1100010000110010: color_data = 12'b001110100111;
		16'b1100010000110011: color_data = 12'b001110100111;
		16'b1100010000110100: color_data = 12'b001110100111;
		16'b1100010000110101: color_data = 12'b001110100111;
		16'b1100010000110110: color_data = 12'b001110100111;
		16'b1100010000110111: color_data = 12'b001110100111;
		16'b1100010001000100: color_data = 12'b001110100111;
		16'b1100010001000101: color_data = 12'b001110100111;
		16'b1100010001000110: color_data = 12'b001110100111;
		16'b1100010001000111: color_data = 12'b001110100111;
		16'b1100010001001000: color_data = 12'b001110100111;
		16'b1100010001001001: color_data = 12'b001110100111;
		16'b1100010001001010: color_data = 12'b001110100111;
		16'b1100010001001011: color_data = 12'b001110100111;
		16'b1100010001001100: color_data = 12'b001110100111;
		16'b1100010001001101: color_data = 12'b001110100111;
		16'b1100010001001110: color_data = 12'b001110100111;
		16'b1100010001001111: color_data = 12'b001110100111;
		16'b1100010001010110: color_data = 12'b001110100111;
		16'b1100010001010111: color_data = 12'b001110100111;
		16'b1100010001011000: color_data = 12'b001110100111;
		16'b1100010001011001: color_data = 12'b001110100111;
		16'b1100010001011010: color_data = 12'b001110100111;
		16'b1100010001011011: color_data = 12'b001110100111;
		16'b1100010001011100: color_data = 12'b001110100111;
		16'b1100010001011101: color_data = 12'b001110100111;
		16'b1100010001011110: color_data = 12'b001110100111;
		16'b1100010001011111: color_data = 12'b001110100111;
		16'b1100010001100000: color_data = 12'b001110100111;
		16'b1100010001100001: color_data = 12'b001110100111;
		16'b1100010001100010: color_data = 12'b001110100111;
		16'b1100010001100011: color_data = 12'b001110100111;
		16'b1100010001100100: color_data = 12'b001110100111;
		16'b1100010001100101: color_data = 12'b001110100111;
		16'b1100010001100110: color_data = 12'b001110100111;
		16'b1100010001100111: color_data = 12'b001110100111;
		16'b1100010001101000: color_data = 12'b001110100111;
		16'b1100010001101001: color_data = 12'b001110100111;
		16'b1100010001101010: color_data = 12'b001110100111;
		16'b1100010001101011: color_data = 12'b001110100111;
		16'b1100010001101100: color_data = 12'b001110100111;
		16'b1100010001101101: color_data = 12'b001110100111;
		16'b1100010001101110: color_data = 12'b001110100111;
		16'b1100010001110101: color_data = 12'b001110100111;
		16'b1100010001110110: color_data = 12'b001110100111;
		16'b1100010001110111: color_data = 12'b001110100111;
		16'b1100010001111000: color_data = 12'b001110100111;
		16'b1100010001111001: color_data = 12'b001110100111;
		16'b1100010001111010: color_data = 12'b001110100111;
		16'b1100010001111011: color_data = 12'b001110100111;
		16'b1100010001111100: color_data = 12'b001110100111;
		16'b1100010001111101: color_data = 12'b001110100111;
		16'b1100010001111110: color_data = 12'b001110100111;
		16'b1100010001111111: color_data = 12'b001110100111;
		16'b1100010010000000: color_data = 12'b001110100111;
		16'b1100010010001101: color_data = 12'b001110100111;
		16'b1100010010001110: color_data = 12'b001110100111;
		16'b1100010010001111: color_data = 12'b001110100111;
		16'b1100010010010000: color_data = 12'b001110100111;
		16'b1100010010010001: color_data = 12'b001110100111;
		16'b1100010010010010: color_data = 12'b001110100111;
		16'b1100010010010011: color_data = 12'b001110100111;
		16'b1100010010010100: color_data = 12'b001110100111;
		16'b1100010010010101: color_data = 12'b001110100111;
		16'b1100010010010110: color_data = 12'b001110100111;
		16'b1100010010010111: color_data = 12'b001110100111;
		16'b1100010010011000: color_data = 12'b001110100111;
		16'b1100010010011001: color_data = 12'b001110100111;
		16'b1100010010100000: color_data = 12'b001110100111;
		16'b1100010010100001: color_data = 12'b001110100111;
		16'b1100010010100010: color_data = 12'b001110100111;
		16'b1100010010100011: color_data = 12'b001110100111;
		16'b1100010010100100: color_data = 12'b001110100111;
		16'b1100010010100101: color_data = 12'b001110100111;
		16'b1100010010100110: color_data = 12'b001110100111;
		16'b1100010010100111: color_data = 12'b001110100111;
		16'b1100010010101000: color_data = 12'b001110100111;
		16'b1100010010101001: color_data = 12'b001110100111;
		16'b1100010010101010: color_data = 12'b001110100111;
		16'b1100010010101011: color_data = 12'b001110100111;
		16'b1100010010101100: color_data = 12'b001110100111;
		16'b1100010010101101: color_data = 12'b001110100111;
		16'b1100010010101110: color_data = 12'b001110100111;
		16'b1100010010101111: color_data = 12'b001110100111;
		16'b1100010010110000: color_data = 12'b001110100111;
		16'b1100010010110001: color_data = 12'b001110100111;
		16'b1100010010110010: color_data = 12'b001110100111;
		16'b1100010010110011: color_data = 12'b001110100111;
		16'b1100010010110100: color_data = 12'b001110100111;
		16'b1100010010110101: color_data = 12'b001110100111;
		16'b1100010010110110: color_data = 12'b001110100111;
		16'b1100010010110111: color_data = 12'b001110100111;
		16'b1100010010111000: color_data = 12'b001110100111;
		16'b1100010010111001: color_data = 12'b001110100111;
		16'b1100010010111010: color_data = 12'b001110100111;
		16'b1100010010111011: color_data = 12'b001110100111;
		16'b1100010010111100: color_data = 12'b001110100111;
		16'b1100010010111101: color_data = 12'b001110100111;
		16'b1100010010111110: color_data = 12'b001110100111;
		16'b1100010010111111: color_data = 12'b001110100111;
		16'b1100010011000000: color_data = 12'b001110100111;
		16'b1100010011000001: color_data = 12'b001110100111;
		16'b1100010011000010: color_data = 12'b001110100111;
		16'b1100010011000011: color_data = 12'b001110100111;
		16'b1100010011000100: color_data = 12'b001110100111;
		16'b1100010011001011: color_data = 12'b001110100111;
		16'b1100010011001100: color_data = 12'b001110100111;
		16'b1100010011001101: color_data = 12'b001110100111;
		16'b1100010011001110: color_data = 12'b001110100111;
		16'b1100010011001111: color_data = 12'b001110100111;
		16'b1100010011010000: color_data = 12'b001110100111;
		16'b1100010011010001: color_data = 12'b001110100111;
		16'b1100010011010010: color_data = 12'b001110100111;
		16'b1100010011010011: color_data = 12'b001110100111;
		16'b1100010011010100: color_data = 12'b001110100111;
		16'b1100010011010101: color_data = 12'b001110100111;
		16'b1100010011010110: color_data = 12'b001110100111;
		16'b1100010011111100: color_data = 12'b001110100111;
		16'b1100010011111101: color_data = 12'b001110100111;
		16'b1100010011111110: color_data = 12'b001110100111;
		16'b1100010011111111: color_data = 12'b001110100111;
		16'b1100010100000000: color_data = 12'b001110100111;
		16'b1100010100000001: color_data = 12'b001110100111;
		16'b1100010100000010: color_data = 12'b001110100111;
		16'b1100010100000011: color_data = 12'b001110100111;
		16'b1100010100000100: color_data = 12'b001110100111;
		16'b1100010100000101: color_data = 12'b001110100111;
		16'b1100010100000110: color_data = 12'b001110100111;
		16'b1100010100000111: color_data = 12'b001110100111;
		16'b1100010100001000: color_data = 12'b001110100111;
		16'b1100010100001001: color_data = 12'b001110100111;
		16'b1100010100001010: color_data = 12'b001110100111;
		16'b1100010100001011: color_data = 12'b001110100111;
		16'b1100010100001100: color_data = 12'b001110100111;
		16'b1100010100001101: color_data = 12'b001110100111;
		16'b1100010100001110: color_data = 12'b001110100111;
		16'b1100010100001111: color_data = 12'b001110100111;
		16'b1100010100010000: color_data = 12'b001110100111;
		16'b1100010100010001: color_data = 12'b001110100111;
		16'b1100010100010010: color_data = 12'b001110100111;
		16'b1100010100010011: color_data = 12'b001110100111;
		16'b1100010100010100: color_data = 12'b001110100111;
		16'b1100010100010101: color_data = 12'b001110100111;
		16'b1100010100010110: color_data = 12'b001110100111;
		16'b1100010100010111: color_data = 12'b001110100111;
		16'b1100010100011000: color_data = 12'b001110100111;
		16'b1100010100011001: color_data = 12'b001110100111;
		16'b1100010100011010: color_data = 12'b001110100111;
		16'b1100010100011011: color_data = 12'b001110100111;
		16'b1100010100011100: color_data = 12'b001110100111;
		16'b1100010100011101: color_data = 12'b001110100111;
		16'b1100010100011110: color_data = 12'b001110100111;
		16'b1100010100011111: color_data = 12'b001110100111;
		16'b1100010100100000: color_data = 12'b001110100111;
		16'b1100010100101101: color_data = 12'b001110100111;
		16'b1100010100101110: color_data = 12'b001110100111;
		16'b1100010100101111: color_data = 12'b001110100111;
		16'b1100010100110000: color_data = 12'b001110100111;
		16'b1100010100110001: color_data = 12'b001110100111;
		16'b1100010100110010: color_data = 12'b001110100111;
		16'b1100010100110011: color_data = 12'b001110100111;
		16'b1100010100110100: color_data = 12'b001110100111;
		16'b1100010100110101: color_data = 12'b001110100111;
		16'b1100010100110110: color_data = 12'b001110100111;
		16'b1100010100110111: color_data = 12'b001110100111;
		16'b1100010100111000: color_data = 12'b001110100111;
		16'b1100010101000101: color_data = 12'b001110100111;
		16'b1100010101000110: color_data = 12'b001110100111;
		16'b1100010101000111: color_data = 12'b001110100111;
		16'b1100010101001000: color_data = 12'b001110100111;
		16'b1100010101001001: color_data = 12'b001110100111;
		16'b1100010101001010: color_data = 12'b001110100111;
		16'b1100010101001011: color_data = 12'b001110100111;
		16'b1100010101001100: color_data = 12'b001110100111;
		16'b1100010101001101: color_data = 12'b001110100111;
		16'b1100010101001110: color_data = 12'b001110100111;
		16'b1100010101001111: color_data = 12'b001110100111;
		16'b1100010101010000: color_data = 12'b001110100111;
		16'b1100010101010001: color_data = 12'b001110100111;
		16'b1100010101011000: color_data = 12'b001110100111;
		16'b1100010101011001: color_data = 12'b001110100111;
		16'b1100010101011010: color_data = 12'b001110100111;
		16'b1100010101011011: color_data = 12'b001110100111;
		16'b1100010101011100: color_data = 12'b001110100111;
		16'b1100010101011101: color_data = 12'b001110100111;
		16'b1100010101011110: color_data = 12'b001110100111;
		16'b1100010101011111: color_data = 12'b001110100111;
		16'b1100010101100000: color_data = 12'b001110100111;
		16'b1100010101100001: color_data = 12'b001110100111;
		16'b1100010101100010: color_data = 12'b001110100111;
		16'b1100010101100011: color_data = 12'b001110100111;
		16'b1100010101100100: color_data = 12'b001110100111;
		16'b1100010101100101: color_data = 12'b001110100111;
		16'b1100010101100110: color_data = 12'b001110100111;
		16'b1100010101100111: color_data = 12'b001110100111;
		16'b1100010101101000: color_data = 12'b001110100111;
		16'b1100010101101001: color_data = 12'b001110100111;
		16'b1100010101101010: color_data = 12'b001110100111;
		16'b1100010101101011: color_data = 12'b001110100111;
		16'b1100010101101100: color_data = 12'b001110100111;
		16'b1100010101101101: color_data = 12'b001110100111;
		16'b1100010101101110: color_data = 12'b001110100111;
		16'b1100010101101111: color_data = 12'b001110100111;
		16'b1100010101110000: color_data = 12'b001110100111;
		16'b1100010101110001: color_data = 12'b001110100111;
		16'b1100010101110010: color_data = 12'b001110100111;
		16'b1100010101110011: color_data = 12'b001110100111;
		16'b1100010101110100: color_data = 12'b001110100111;
		16'b1100010101110101: color_data = 12'b001110100111;
		16'b1100010101110110: color_data = 12'b001110100111;
		16'b1100010101110111: color_data = 12'b001110100111;
		16'b1100010101111000: color_data = 12'b001110100111;
		16'b1100010101111001: color_data = 12'b001110100111;
		16'b1100010101111010: color_data = 12'b001110100111;
		16'b1100010101111011: color_data = 12'b001110100111;
		16'b1100011000000000: color_data = 12'b001110100111;
		16'b1100011000000001: color_data = 12'b001110100111;
		16'b1100011000000010: color_data = 12'b001110100111;
		16'b1100011000000011: color_data = 12'b001110100111;
		16'b1100011000000100: color_data = 12'b001110100111;
		16'b1100011000000101: color_data = 12'b001110100111;
		16'b1100011000000110: color_data = 12'b001110100111;
		16'b1100011000000111: color_data = 12'b001110100111;
		16'b1100011000001000: color_data = 12'b001110100111;
		16'b1100011000001001: color_data = 12'b001110100111;
		16'b1100011000001010: color_data = 12'b001110100111;
		16'b1100011000001011: color_data = 12'b001110100111;
		16'b1100011000001100: color_data = 12'b001110100111;
		16'b1100011000001101: color_data = 12'b001110100111;
		16'b1100011000001110: color_data = 12'b001110100111;
		16'b1100011000001111: color_data = 12'b001110100111;
		16'b1100011000010000: color_data = 12'b001110100111;
		16'b1100011000010001: color_data = 12'b001110100111;
		16'b1100011000010010: color_data = 12'b001110100111;
		16'b1100011000010011: color_data = 12'b001110100111;
		16'b1100011000010100: color_data = 12'b001110100111;
		16'b1100011000010101: color_data = 12'b001110100111;
		16'b1100011000010110: color_data = 12'b001110100111;
		16'b1100011000010111: color_data = 12'b001110100111;
		16'b1100011000011000: color_data = 12'b001110100111;
		16'b1100011000011001: color_data = 12'b001110100111;
		16'b1100011000011010: color_data = 12'b001110100111;
		16'b1100011000011011: color_data = 12'b001110100111;
		16'b1100011000011100: color_data = 12'b001110100111;
		16'b1100011000011101: color_data = 12'b001110100111;
		16'b1100011000011110: color_data = 12'b001110100111;
		16'b1100011000011111: color_data = 12'b001110100111;
		16'b1100011000100000: color_data = 12'b001110100111;
		16'b1100011000100001: color_data = 12'b001110100111;
		16'b1100011000100010: color_data = 12'b001110100111;
		16'b1100011000100011: color_data = 12'b001110100111;
		16'b1100011000100100: color_data = 12'b001110100111;
		16'b1100011000101011: color_data = 12'b001110100111;
		16'b1100011000101100: color_data = 12'b001110100111;
		16'b1100011000101101: color_data = 12'b001110100111;
		16'b1100011000101110: color_data = 12'b001110100111;
		16'b1100011000101111: color_data = 12'b001110100111;
		16'b1100011000110000: color_data = 12'b001110100111;
		16'b1100011000110001: color_data = 12'b001110100111;
		16'b1100011000110010: color_data = 12'b001110100111;
		16'b1100011000110011: color_data = 12'b001110100111;
		16'b1100011000110100: color_data = 12'b001110100111;
		16'b1100011000110101: color_data = 12'b001110100111;
		16'b1100011000110110: color_data = 12'b001110100111;
		16'b1100011000110111: color_data = 12'b001110100111;
		16'b1100011001000100: color_data = 12'b001110100111;
		16'b1100011001000101: color_data = 12'b001110100111;
		16'b1100011001000110: color_data = 12'b001110100111;
		16'b1100011001000111: color_data = 12'b001110100111;
		16'b1100011001001000: color_data = 12'b001110100111;
		16'b1100011001001001: color_data = 12'b001110100111;
		16'b1100011001001010: color_data = 12'b001110100111;
		16'b1100011001001011: color_data = 12'b001110100111;
		16'b1100011001001100: color_data = 12'b001110100111;
		16'b1100011001001101: color_data = 12'b001110100111;
		16'b1100011001001110: color_data = 12'b001110100111;
		16'b1100011001001111: color_data = 12'b001110100111;
		16'b1100011001010110: color_data = 12'b001110100111;
		16'b1100011001010111: color_data = 12'b001110100111;
		16'b1100011001011000: color_data = 12'b001110100111;
		16'b1100011001011001: color_data = 12'b001110100111;
		16'b1100011001011010: color_data = 12'b001110100111;
		16'b1100011001011011: color_data = 12'b001110100111;
		16'b1100011001011100: color_data = 12'b001110100111;
		16'b1100011001011101: color_data = 12'b001110100111;
		16'b1100011001011110: color_data = 12'b001110100111;
		16'b1100011001011111: color_data = 12'b001110100111;
		16'b1100011001100000: color_data = 12'b001110100111;
		16'b1100011001100001: color_data = 12'b001110100111;
		16'b1100011001100010: color_data = 12'b001110100111;
		16'b1100011001100011: color_data = 12'b001110100111;
		16'b1100011001100100: color_data = 12'b001110100111;
		16'b1100011001100101: color_data = 12'b001110100111;
		16'b1100011001100110: color_data = 12'b001110100111;
		16'b1100011001100111: color_data = 12'b001110100111;
		16'b1100011001101000: color_data = 12'b001110100111;
		16'b1100011001101001: color_data = 12'b001110100111;
		16'b1100011001101010: color_data = 12'b001110100111;
		16'b1100011001101011: color_data = 12'b001110100111;
		16'b1100011001101100: color_data = 12'b001110100111;
		16'b1100011001101101: color_data = 12'b001110100111;
		16'b1100011001101110: color_data = 12'b001110100111;
		16'b1100011001110101: color_data = 12'b001110100111;
		16'b1100011001110110: color_data = 12'b001110100111;
		16'b1100011001110111: color_data = 12'b001110100111;
		16'b1100011001111000: color_data = 12'b001110100111;
		16'b1100011001111001: color_data = 12'b001110100111;
		16'b1100011001111010: color_data = 12'b001110100111;
		16'b1100011001111011: color_data = 12'b001110100111;
		16'b1100011001111100: color_data = 12'b001110100111;
		16'b1100011001111101: color_data = 12'b001110100111;
		16'b1100011001111110: color_data = 12'b001110100111;
		16'b1100011001111111: color_data = 12'b001110100111;
		16'b1100011010000000: color_data = 12'b001110100111;
		16'b1100011010001101: color_data = 12'b001110100111;
		16'b1100011010001110: color_data = 12'b001110100111;
		16'b1100011010001111: color_data = 12'b001110100111;
		16'b1100011010010000: color_data = 12'b001110100111;
		16'b1100011010010001: color_data = 12'b001110100111;
		16'b1100011010010010: color_data = 12'b001110100111;
		16'b1100011010010011: color_data = 12'b001110100111;
		16'b1100011010010100: color_data = 12'b001110100111;
		16'b1100011010010101: color_data = 12'b001110100111;
		16'b1100011010010110: color_data = 12'b001110100111;
		16'b1100011010010111: color_data = 12'b001110100111;
		16'b1100011010011000: color_data = 12'b001110100111;
		16'b1100011010011001: color_data = 12'b001110100111;
		16'b1100011010100000: color_data = 12'b001110100111;
		16'b1100011010100001: color_data = 12'b001110100111;
		16'b1100011010100010: color_data = 12'b001110100111;
		16'b1100011010100011: color_data = 12'b001110100111;
		16'b1100011010100100: color_data = 12'b001110100111;
		16'b1100011010100101: color_data = 12'b001110100111;
		16'b1100011010100110: color_data = 12'b001110100111;
		16'b1100011010100111: color_data = 12'b001110100111;
		16'b1100011010101000: color_data = 12'b001110100111;
		16'b1100011010101001: color_data = 12'b001110100111;
		16'b1100011010101010: color_data = 12'b001110100111;
		16'b1100011010101011: color_data = 12'b001110100111;
		16'b1100011010101100: color_data = 12'b001110100111;
		16'b1100011010101101: color_data = 12'b001110100111;
		16'b1100011010101110: color_data = 12'b001110100111;
		16'b1100011010101111: color_data = 12'b001110100111;
		16'b1100011010110000: color_data = 12'b001110100111;
		16'b1100011010110001: color_data = 12'b001110100111;
		16'b1100011010110010: color_data = 12'b001110100111;
		16'b1100011010110011: color_data = 12'b001110100111;
		16'b1100011010110100: color_data = 12'b001110100111;
		16'b1100011010110101: color_data = 12'b001110100111;
		16'b1100011010110110: color_data = 12'b001110100111;
		16'b1100011010110111: color_data = 12'b001110100111;
		16'b1100011010111000: color_data = 12'b001110100111;
		16'b1100011010111001: color_data = 12'b001110100111;
		16'b1100011010111010: color_data = 12'b001110100111;
		16'b1100011010111011: color_data = 12'b001110100111;
		16'b1100011010111100: color_data = 12'b001110100111;
		16'b1100011010111101: color_data = 12'b001110100111;
		16'b1100011010111110: color_data = 12'b001110100111;
		16'b1100011010111111: color_data = 12'b001110100111;
		16'b1100011011000000: color_data = 12'b001110100111;
		16'b1100011011000001: color_data = 12'b001110100111;
		16'b1100011011000010: color_data = 12'b001110100111;
		16'b1100011011000011: color_data = 12'b001110100111;
		16'b1100011011000100: color_data = 12'b001110100111;
		16'b1100011011001011: color_data = 12'b001110100111;
		16'b1100011011001100: color_data = 12'b001110100111;
		16'b1100011011001101: color_data = 12'b001110100111;
		16'b1100011011001110: color_data = 12'b001110100111;
		16'b1100011011001111: color_data = 12'b001110100111;
		16'b1100011011010000: color_data = 12'b001110100111;
		16'b1100011011010001: color_data = 12'b001110100111;
		16'b1100011011010010: color_data = 12'b001110100111;
		16'b1100011011010011: color_data = 12'b001110100111;
		16'b1100011011010100: color_data = 12'b001110100111;
		16'b1100011011010101: color_data = 12'b001110100111;
		16'b1100011011010110: color_data = 12'b001110100111;
		16'b1100011011111100: color_data = 12'b001110100111;
		16'b1100011011111101: color_data = 12'b001110100111;
		16'b1100011011111110: color_data = 12'b001110100111;
		16'b1100011011111111: color_data = 12'b001110100111;
		16'b1100011100000000: color_data = 12'b001110100111;
		16'b1100011100000001: color_data = 12'b001110100111;
		16'b1100011100000010: color_data = 12'b001110100111;
		16'b1100011100000011: color_data = 12'b001110100111;
		16'b1100011100000100: color_data = 12'b001110100111;
		16'b1100011100000101: color_data = 12'b001110100111;
		16'b1100011100000110: color_data = 12'b001110100111;
		16'b1100011100000111: color_data = 12'b001110100111;
		16'b1100011100001000: color_data = 12'b001110100111;
		16'b1100011100001001: color_data = 12'b001110100111;
		16'b1100011100001010: color_data = 12'b001110100111;
		16'b1100011100001011: color_data = 12'b001110100111;
		16'b1100011100001100: color_data = 12'b001110100111;
		16'b1100011100001101: color_data = 12'b001110100111;
		16'b1100011100001110: color_data = 12'b001110100111;
		16'b1100011100001111: color_data = 12'b001110100111;
		16'b1100011100010000: color_data = 12'b001110100111;
		16'b1100011100010001: color_data = 12'b001110100111;
		16'b1100011100010010: color_data = 12'b001110100111;
		16'b1100011100010011: color_data = 12'b001110100111;
		16'b1100011100010100: color_data = 12'b001110100111;
		16'b1100011100010101: color_data = 12'b001110100111;
		16'b1100011100010110: color_data = 12'b001110100111;
		16'b1100011100010111: color_data = 12'b001110100111;
		16'b1100011100011000: color_data = 12'b001110100111;
		16'b1100011100011001: color_data = 12'b001110100111;
		16'b1100011100011010: color_data = 12'b001110100111;
		16'b1100011100011011: color_data = 12'b001110100111;
		16'b1100011100011100: color_data = 12'b001110100111;
		16'b1100011100011101: color_data = 12'b001110100111;
		16'b1100011100011110: color_data = 12'b001110100111;
		16'b1100011100011111: color_data = 12'b001110100111;
		16'b1100011100100000: color_data = 12'b001110100111;
		16'b1100011100101101: color_data = 12'b001110100111;
		16'b1100011100101110: color_data = 12'b001110100111;
		16'b1100011100101111: color_data = 12'b001110100111;
		16'b1100011100110000: color_data = 12'b001110100111;
		16'b1100011100110001: color_data = 12'b001110100111;
		16'b1100011100110010: color_data = 12'b001110100111;
		16'b1100011100110011: color_data = 12'b001110100111;
		16'b1100011100110100: color_data = 12'b001110100111;
		16'b1100011100110101: color_data = 12'b001110100111;
		16'b1100011100110110: color_data = 12'b001110100111;
		16'b1100011100110111: color_data = 12'b001110100111;
		16'b1100011100111000: color_data = 12'b001110100111;
		16'b1100011101000101: color_data = 12'b001110100111;
		16'b1100011101000110: color_data = 12'b001110100111;
		16'b1100011101000111: color_data = 12'b001110100111;
		16'b1100011101001000: color_data = 12'b001110100111;
		16'b1100011101001001: color_data = 12'b001110100111;
		16'b1100011101001010: color_data = 12'b001110100111;
		16'b1100011101001011: color_data = 12'b001110100111;
		16'b1100011101001100: color_data = 12'b001110100111;
		16'b1100011101001101: color_data = 12'b001110100111;
		16'b1100011101001110: color_data = 12'b001110100111;
		16'b1100011101001111: color_data = 12'b001110100111;
		16'b1100011101010000: color_data = 12'b001110100111;
		16'b1100011101010001: color_data = 12'b001110100111;
		16'b1100011101011000: color_data = 12'b001110100111;
		16'b1100011101011001: color_data = 12'b001110100111;
		16'b1100011101011010: color_data = 12'b001110100111;
		16'b1100011101011011: color_data = 12'b001110100111;
		16'b1100011101011100: color_data = 12'b001110100111;
		16'b1100011101011101: color_data = 12'b001110100111;
		16'b1100011101011110: color_data = 12'b001110100111;
		16'b1100011101011111: color_data = 12'b001110100111;
		16'b1100011101100000: color_data = 12'b001110100111;
		16'b1100011101100001: color_data = 12'b001110100111;
		16'b1100011101100010: color_data = 12'b001110100111;
		16'b1100011101100011: color_data = 12'b001110100111;
		16'b1100011101100100: color_data = 12'b001110100111;
		16'b1100011101100101: color_data = 12'b001110100111;
		16'b1100011101100110: color_data = 12'b001110100111;
		16'b1100011101100111: color_data = 12'b001110100111;
		16'b1100011101101000: color_data = 12'b001110100111;
		16'b1100011101101001: color_data = 12'b001110100111;
		16'b1100011101101010: color_data = 12'b001110100111;
		16'b1100011101101011: color_data = 12'b001110100111;
		16'b1100011101101100: color_data = 12'b001110100111;
		16'b1100011101101101: color_data = 12'b001110100111;
		16'b1100011101101110: color_data = 12'b001110100111;
		16'b1100011101101111: color_data = 12'b001110100111;
		16'b1100011101110000: color_data = 12'b001110100111;
		16'b1100011101110001: color_data = 12'b001110100111;
		16'b1100011101110010: color_data = 12'b001110100111;
		16'b1100011101110011: color_data = 12'b001110100111;
		16'b1100011101110100: color_data = 12'b001110100111;
		16'b1100011101110101: color_data = 12'b001110100111;
		16'b1100011101110110: color_data = 12'b001110100111;
		16'b1100011101110111: color_data = 12'b001110100111;
		16'b1100011101111000: color_data = 12'b001110100111;
		16'b1100011101111001: color_data = 12'b001110100111;
		16'b1100011101111010: color_data = 12'b001110100111;
		16'b1100011101111011: color_data = 12'b001110100111;
		16'b1100100000000000: color_data = 12'b001110100111;
		16'b1100100000000001: color_data = 12'b001110100111;
		16'b1100100000000010: color_data = 12'b001110100111;
		16'b1100100000000011: color_data = 12'b001110100111;
		16'b1100100000000100: color_data = 12'b001110100111;
		16'b1100100000000101: color_data = 12'b001110100111;
		16'b1100100000000110: color_data = 12'b001110100111;
		16'b1100100000000111: color_data = 12'b001110100111;
		16'b1100100000001000: color_data = 12'b001110100111;
		16'b1100100000001001: color_data = 12'b001110100111;
		16'b1100100000001010: color_data = 12'b001110100111;
		16'b1100100000001011: color_data = 12'b001110100111;
		16'b1100100000001100: color_data = 12'b001110100111;
		16'b1100100000001101: color_data = 12'b001110100111;
		16'b1100100000001110: color_data = 12'b001110100111;
		16'b1100100000001111: color_data = 12'b001110100111;
		16'b1100100000010000: color_data = 12'b001110100111;
		16'b1100100000010001: color_data = 12'b001110100111;
		16'b1100100000010010: color_data = 12'b001110100111;
		16'b1100100000010011: color_data = 12'b001110100111;
		16'b1100100000010100: color_data = 12'b001110100111;
		16'b1100100000010101: color_data = 12'b001110100111;
		16'b1100100000010110: color_data = 12'b001110100111;
		16'b1100100000010111: color_data = 12'b001110100111;
		16'b1100100000011000: color_data = 12'b001110100111;
		16'b1100100000011001: color_data = 12'b001110100111;
		16'b1100100000011010: color_data = 12'b001110100111;
		16'b1100100000011011: color_data = 12'b001110100111;
		16'b1100100000011100: color_data = 12'b001110100111;
		16'b1100100000011101: color_data = 12'b001110100111;
		16'b1100100000011110: color_data = 12'b001110100111;
		16'b1100100000011111: color_data = 12'b001110100111;
		16'b1100100000100000: color_data = 12'b001110100111;
		16'b1100100000100001: color_data = 12'b001110100111;
		16'b1100100000100010: color_data = 12'b001110100111;
		16'b1100100000100011: color_data = 12'b001110100111;
		16'b1100100000100100: color_data = 12'b001110100111;
		16'b1100100000101011: color_data = 12'b001110100111;
		16'b1100100000101100: color_data = 12'b001110100111;
		16'b1100100000101101: color_data = 12'b001110100111;
		16'b1100100000101110: color_data = 12'b001110100111;
		16'b1100100000101111: color_data = 12'b001110100111;
		16'b1100100000110000: color_data = 12'b001110100111;
		16'b1100100000110001: color_data = 12'b001110100111;
		16'b1100100000110010: color_data = 12'b001110100111;
		16'b1100100000110011: color_data = 12'b001110100111;
		16'b1100100000110100: color_data = 12'b001110100111;
		16'b1100100000110101: color_data = 12'b001110100111;
		16'b1100100000110110: color_data = 12'b001110100111;
		16'b1100100000110111: color_data = 12'b001110100111;
		16'b1100100001000100: color_data = 12'b001110100111;
		16'b1100100001000101: color_data = 12'b001110100111;
		16'b1100100001000110: color_data = 12'b001110100111;
		16'b1100100001000111: color_data = 12'b001110100111;
		16'b1100100001001000: color_data = 12'b001110100111;
		16'b1100100001001001: color_data = 12'b001110100111;
		16'b1100100001001010: color_data = 12'b001110100111;
		16'b1100100001001011: color_data = 12'b001110100111;
		16'b1100100001001100: color_data = 12'b001110100111;
		16'b1100100001001101: color_data = 12'b001110100111;
		16'b1100100001001110: color_data = 12'b001110100111;
		16'b1100100001001111: color_data = 12'b001110100111;
		16'b1100100001010110: color_data = 12'b001110100111;
		16'b1100100001010111: color_data = 12'b001110100111;
		16'b1100100001011000: color_data = 12'b001110100111;
		16'b1100100001011001: color_data = 12'b001110100111;
		16'b1100100001011010: color_data = 12'b001110100111;
		16'b1100100001011011: color_data = 12'b001110100111;
		16'b1100100001011100: color_data = 12'b001110100111;
		16'b1100100001011101: color_data = 12'b001110100111;
		16'b1100100001011110: color_data = 12'b001110100111;
		16'b1100100001011111: color_data = 12'b001110100111;
		16'b1100100001100000: color_data = 12'b001110100111;
		16'b1100100001100001: color_data = 12'b001110100111;
		16'b1100100001100010: color_data = 12'b001110100111;
		16'b1100100001100011: color_data = 12'b001110100111;
		16'b1100100001100100: color_data = 12'b001110100111;
		16'b1100100001100101: color_data = 12'b001110100111;
		16'b1100100001100110: color_data = 12'b001110100111;
		16'b1100100001100111: color_data = 12'b001110100111;
		16'b1100100001101000: color_data = 12'b001110100111;
		16'b1100100001101001: color_data = 12'b001110100111;
		16'b1100100001101010: color_data = 12'b001110100111;
		16'b1100100001101011: color_data = 12'b001110100111;
		16'b1100100001101100: color_data = 12'b001110100111;
		16'b1100100001101101: color_data = 12'b001110100111;
		16'b1100100001101110: color_data = 12'b001110100111;
		16'b1100100001110101: color_data = 12'b001110100111;
		16'b1100100001110110: color_data = 12'b001110100111;
		16'b1100100001110111: color_data = 12'b001110100111;
		16'b1100100001111000: color_data = 12'b001110100111;
		16'b1100100001111001: color_data = 12'b001110100111;
		16'b1100100001111010: color_data = 12'b001110100111;
		16'b1100100001111011: color_data = 12'b001110100111;
		16'b1100100001111100: color_data = 12'b001110100111;
		16'b1100100001111101: color_data = 12'b001110100111;
		16'b1100100001111110: color_data = 12'b001110100111;
		16'b1100100001111111: color_data = 12'b001110100111;
		16'b1100100010000000: color_data = 12'b001110100111;
		16'b1100100010001101: color_data = 12'b001110100111;
		16'b1100100010001110: color_data = 12'b001110100111;
		16'b1100100010001111: color_data = 12'b001110100111;
		16'b1100100010010000: color_data = 12'b001110100111;
		16'b1100100010010001: color_data = 12'b001110100111;
		16'b1100100010010010: color_data = 12'b001110100111;
		16'b1100100010010011: color_data = 12'b001110100111;
		16'b1100100010010100: color_data = 12'b001110100111;
		16'b1100100010010101: color_data = 12'b001110100111;
		16'b1100100010010110: color_data = 12'b001110100111;
		16'b1100100010010111: color_data = 12'b001110100111;
		16'b1100100010011000: color_data = 12'b001110100111;
		16'b1100100010011001: color_data = 12'b001110100111;
		16'b1100100010100000: color_data = 12'b001110100111;
		16'b1100100010100001: color_data = 12'b001110100111;
		16'b1100100010100010: color_data = 12'b001110100111;
		16'b1100100010100011: color_data = 12'b001110100111;
		16'b1100100010100100: color_data = 12'b001110100111;
		16'b1100100010100101: color_data = 12'b001110100111;
		16'b1100100010100110: color_data = 12'b001110100111;
		16'b1100100010100111: color_data = 12'b001110100111;
		16'b1100100010101000: color_data = 12'b001110100111;
		16'b1100100010101001: color_data = 12'b001110100111;
		16'b1100100010101010: color_data = 12'b001110100111;
		16'b1100100010101011: color_data = 12'b001110100111;
		16'b1100100010101100: color_data = 12'b001110100111;
		16'b1100100010101101: color_data = 12'b001110100111;
		16'b1100100010101110: color_data = 12'b001110100111;
		16'b1100100010101111: color_data = 12'b001110100111;
		16'b1100100010110000: color_data = 12'b001110100111;
		16'b1100100010110001: color_data = 12'b001110100111;
		16'b1100100010110010: color_data = 12'b001110100111;
		16'b1100100010110011: color_data = 12'b001110100111;
		16'b1100100010110100: color_data = 12'b001110100111;
		16'b1100100010110101: color_data = 12'b001110100111;
		16'b1100100010110110: color_data = 12'b001110100111;
		16'b1100100010110111: color_data = 12'b001110100111;
		16'b1100100010111000: color_data = 12'b001110100111;
		16'b1100100010111001: color_data = 12'b001110100111;
		16'b1100100010111010: color_data = 12'b001110100111;
		16'b1100100010111011: color_data = 12'b001110100111;
		16'b1100100010111100: color_data = 12'b001110100111;
		16'b1100100010111101: color_data = 12'b001110100111;
		16'b1100100010111110: color_data = 12'b001110100111;
		16'b1100100010111111: color_data = 12'b001110100111;
		16'b1100100011000000: color_data = 12'b001110100111;
		16'b1100100011000001: color_data = 12'b001110100111;
		16'b1100100011000010: color_data = 12'b001110100111;
		16'b1100100011000011: color_data = 12'b001110100111;
		16'b1100100011000100: color_data = 12'b001110100111;
		16'b1100100011001011: color_data = 12'b001110100111;
		16'b1100100011001100: color_data = 12'b001110100111;
		16'b1100100011001101: color_data = 12'b001110100111;
		16'b1100100011001110: color_data = 12'b001110100111;
		16'b1100100011001111: color_data = 12'b001110100111;
		16'b1100100011010000: color_data = 12'b001110100111;
		16'b1100100011010001: color_data = 12'b001110100111;
		16'b1100100011010010: color_data = 12'b001110100111;
		16'b1100100011010011: color_data = 12'b001110100111;
		16'b1100100011010100: color_data = 12'b001110100111;
		16'b1100100011010101: color_data = 12'b001110100111;
		16'b1100100011010110: color_data = 12'b001110100111;
		16'b1100100011111100: color_data = 12'b001110100111;
		16'b1100100011111101: color_data = 12'b001110100111;
		16'b1100100011111110: color_data = 12'b001110100111;
		16'b1100100011111111: color_data = 12'b001110100111;
		16'b1100100100000000: color_data = 12'b001110100111;
		16'b1100100100000001: color_data = 12'b001110100111;
		16'b1100100100000010: color_data = 12'b001110100111;
		16'b1100100100000011: color_data = 12'b001110100111;
		16'b1100100100000100: color_data = 12'b001110100111;
		16'b1100100100000101: color_data = 12'b001110100111;
		16'b1100100100000110: color_data = 12'b001110100111;
		16'b1100100100000111: color_data = 12'b001110100111;
		16'b1100100100001000: color_data = 12'b001110100111;
		16'b1100100100001001: color_data = 12'b001110100111;
		16'b1100100100001010: color_data = 12'b001110100111;
		16'b1100100100001011: color_data = 12'b001110100111;
		16'b1100100100001100: color_data = 12'b001110100111;
		16'b1100100100001101: color_data = 12'b001110100111;
		16'b1100100100001110: color_data = 12'b001110100111;
		16'b1100100100001111: color_data = 12'b001110100111;
		16'b1100100100010000: color_data = 12'b001110100111;
		16'b1100100100010001: color_data = 12'b001110100111;
		16'b1100100100010010: color_data = 12'b001110100111;
		16'b1100100100010011: color_data = 12'b001110100111;
		16'b1100100100010100: color_data = 12'b001110100111;
		16'b1100100100010101: color_data = 12'b001110100111;
		16'b1100100100010110: color_data = 12'b001110100111;
		16'b1100100100010111: color_data = 12'b001110100111;
		16'b1100100100011000: color_data = 12'b001110100111;
		16'b1100100100011001: color_data = 12'b001110100111;
		16'b1100100100011010: color_data = 12'b001110100111;
		16'b1100100100011011: color_data = 12'b001110100111;
		16'b1100100100011100: color_data = 12'b001110100111;
		16'b1100100100011101: color_data = 12'b001110100111;
		16'b1100100100011110: color_data = 12'b001110100111;
		16'b1100100100011111: color_data = 12'b001110100111;
		16'b1100100100100000: color_data = 12'b001110100111;
		16'b1100100100101101: color_data = 12'b001110100111;
		16'b1100100100101110: color_data = 12'b001110100111;
		16'b1100100100101111: color_data = 12'b001110100111;
		16'b1100100100110000: color_data = 12'b001110100111;
		16'b1100100100110001: color_data = 12'b001110100111;
		16'b1100100100110010: color_data = 12'b001110100111;
		16'b1100100100110011: color_data = 12'b001110100111;
		16'b1100100100110100: color_data = 12'b001110100111;
		16'b1100100100110101: color_data = 12'b001110100111;
		16'b1100100100110110: color_data = 12'b001110100111;
		16'b1100100100110111: color_data = 12'b001110100111;
		16'b1100100100111000: color_data = 12'b001110100111;
		16'b1100100101000101: color_data = 12'b001110100111;
		16'b1100100101000110: color_data = 12'b001110100111;
		16'b1100100101000111: color_data = 12'b001110100111;
		16'b1100100101001000: color_data = 12'b001110100111;
		16'b1100100101001001: color_data = 12'b001110100111;
		16'b1100100101001010: color_data = 12'b001110100111;
		16'b1100100101001011: color_data = 12'b001110100111;
		16'b1100100101001100: color_data = 12'b001110100111;
		16'b1100100101001101: color_data = 12'b001110100111;
		16'b1100100101001110: color_data = 12'b001110100111;
		16'b1100100101001111: color_data = 12'b001110100111;
		16'b1100100101010000: color_data = 12'b001110100111;
		16'b1100100101010001: color_data = 12'b001110100111;
		16'b1100100101011000: color_data = 12'b001110100111;
		16'b1100100101011001: color_data = 12'b001110100111;
		16'b1100100101011010: color_data = 12'b001110100111;
		16'b1100100101011011: color_data = 12'b001110100111;
		16'b1100100101011100: color_data = 12'b001110100111;
		16'b1100100101011101: color_data = 12'b001110100111;
		16'b1100100101011110: color_data = 12'b001110100111;
		16'b1100100101011111: color_data = 12'b001110100111;
		16'b1100100101100000: color_data = 12'b001110100111;
		16'b1100100101100001: color_data = 12'b001110100111;
		16'b1100100101100010: color_data = 12'b001110100111;
		16'b1100100101100011: color_data = 12'b001110100111;
		16'b1100100101100100: color_data = 12'b001110100111;
		16'b1100100101100101: color_data = 12'b001110100111;
		16'b1100100101100110: color_data = 12'b001110100111;
		16'b1100100101100111: color_data = 12'b001110100111;
		16'b1100100101101000: color_data = 12'b001110100111;
		16'b1100100101101001: color_data = 12'b001110100111;
		16'b1100100101101010: color_data = 12'b001110100111;
		16'b1100100101101011: color_data = 12'b001110100111;
		16'b1100100101101100: color_data = 12'b001110100111;
		16'b1100100101101101: color_data = 12'b001110100111;
		16'b1100100101101110: color_data = 12'b001110100111;
		16'b1100100101101111: color_data = 12'b001110100111;
		16'b1100100101110000: color_data = 12'b001110100111;
		16'b1100100101110001: color_data = 12'b001110100111;
		16'b1100100101110010: color_data = 12'b001110100111;
		16'b1100100101110011: color_data = 12'b001110100111;
		16'b1100100101110100: color_data = 12'b001110100111;
		16'b1100100101110101: color_data = 12'b001110100111;
		16'b1100100101110110: color_data = 12'b001110100111;
		16'b1100100101110111: color_data = 12'b001110100111;
		16'b1100100101111000: color_data = 12'b001110100111;
		16'b1100100101111001: color_data = 12'b001110100111;
		16'b1100100101111010: color_data = 12'b001110100111;
		16'b1100100101111011: color_data = 12'b001110100111;
		16'b1100101000000000: color_data = 12'b001110100111;
		16'b1100101000000001: color_data = 12'b001110100111;
		16'b1100101000000010: color_data = 12'b001110100111;
		16'b1100101000000011: color_data = 12'b001110100111;
		16'b1100101000000100: color_data = 12'b001110100111;
		16'b1100101000000101: color_data = 12'b001110100111;
		16'b1100101000000110: color_data = 12'b001110100111;
		16'b1100101000000111: color_data = 12'b001110100111;
		16'b1100101000001000: color_data = 12'b001110100111;
		16'b1100101000001001: color_data = 12'b001110100111;
		16'b1100101000001010: color_data = 12'b001110100111;
		16'b1100101000001011: color_data = 12'b001110100111;
		16'b1100101000001100: color_data = 12'b001110100111;
		16'b1100101000001101: color_data = 12'b001110100111;
		16'b1100101000001110: color_data = 12'b001110100111;
		16'b1100101000001111: color_data = 12'b001110100111;
		16'b1100101000010000: color_data = 12'b001110100111;
		16'b1100101000010001: color_data = 12'b001110100111;
		16'b1100101000010010: color_data = 12'b001110100111;
		16'b1100101000010011: color_data = 12'b001110100111;
		16'b1100101000010100: color_data = 12'b001110100111;
		16'b1100101000010101: color_data = 12'b001110100111;
		16'b1100101000010110: color_data = 12'b001110100111;
		16'b1100101000010111: color_data = 12'b001110100111;
		16'b1100101000011000: color_data = 12'b001110100111;
		16'b1100101000011001: color_data = 12'b001110100111;
		16'b1100101000011010: color_data = 12'b001110100111;
		16'b1100101000011011: color_data = 12'b001110100111;
		16'b1100101000011100: color_data = 12'b001110100111;
		16'b1100101000011101: color_data = 12'b001110100111;
		16'b1100101000011110: color_data = 12'b001110100111;
		16'b1100101000011111: color_data = 12'b001110100111;
		16'b1100101000100000: color_data = 12'b001110100111;
		16'b1100101000100001: color_data = 12'b001110100111;
		16'b1100101000100010: color_data = 12'b001110100111;
		16'b1100101000100011: color_data = 12'b001110100111;
		16'b1100101000100100: color_data = 12'b001110100111;
		16'b1100101000101011: color_data = 12'b001110100111;
		16'b1100101000101100: color_data = 12'b001110100111;
		16'b1100101000101101: color_data = 12'b001110100111;
		16'b1100101000101110: color_data = 12'b001110100111;
		16'b1100101000101111: color_data = 12'b001110100111;
		16'b1100101000110000: color_data = 12'b001110100111;
		16'b1100101000110001: color_data = 12'b001110100111;
		16'b1100101000110010: color_data = 12'b001110100111;
		16'b1100101000110011: color_data = 12'b001110100111;
		16'b1100101000110100: color_data = 12'b001110100111;
		16'b1100101000110101: color_data = 12'b001110100111;
		16'b1100101000110110: color_data = 12'b001110100111;
		16'b1100101000110111: color_data = 12'b001110100111;
		16'b1100101001000100: color_data = 12'b001110100111;
		16'b1100101001000101: color_data = 12'b001110100111;
		16'b1100101001000110: color_data = 12'b001110100111;
		16'b1100101001000111: color_data = 12'b001110100111;
		16'b1100101001001000: color_data = 12'b001110100111;
		16'b1100101001001001: color_data = 12'b001110100111;
		16'b1100101001001010: color_data = 12'b001110100111;
		16'b1100101001001011: color_data = 12'b001110100111;
		16'b1100101001001100: color_data = 12'b001110100111;
		16'b1100101001001101: color_data = 12'b001110100111;
		16'b1100101001001110: color_data = 12'b001110100111;
		16'b1100101001001111: color_data = 12'b001110100111;
		16'b1100101001010110: color_data = 12'b001110100111;
		16'b1100101001010111: color_data = 12'b001110100111;
		16'b1100101001011000: color_data = 12'b001110100111;
		16'b1100101001011001: color_data = 12'b001110100111;
		16'b1100101001011010: color_data = 12'b001110100111;
		16'b1100101001011011: color_data = 12'b001110100111;
		16'b1100101001011100: color_data = 12'b001110100111;
		16'b1100101001011101: color_data = 12'b001110100111;
		16'b1100101001011110: color_data = 12'b001110100111;
		16'b1100101001011111: color_data = 12'b001110100111;
		16'b1100101001100000: color_data = 12'b001110100111;
		16'b1100101001100001: color_data = 12'b001110100111;
		16'b1100101001100010: color_data = 12'b001110100111;
		16'b1100101001100011: color_data = 12'b001110100111;
		16'b1100101001100100: color_data = 12'b001110100111;
		16'b1100101001100101: color_data = 12'b001110100111;
		16'b1100101001100110: color_data = 12'b001110100111;
		16'b1100101001100111: color_data = 12'b001110100111;
		16'b1100101001101000: color_data = 12'b001110100111;
		16'b1100101001101001: color_data = 12'b001110100111;
		16'b1100101001101010: color_data = 12'b001110100111;
		16'b1100101001101011: color_data = 12'b001110100111;
		16'b1100101001101100: color_data = 12'b001110100111;
		16'b1100101001101101: color_data = 12'b001110100111;
		16'b1100101001101110: color_data = 12'b001110100111;
		16'b1100101001110101: color_data = 12'b001110100111;
		16'b1100101001110110: color_data = 12'b001110100111;
		16'b1100101001110111: color_data = 12'b001110100111;
		16'b1100101001111000: color_data = 12'b001110100111;
		16'b1100101001111001: color_data = 12'b001110100111;
		16'b1100101001111010: color_data = 12'b001110100111;
		16'b1100101001111011: color_data = 12'b001110100111;
		16'b1100101001111100: color_data = 12'b001110100111;
		16'b1100101001111101: color_data = 12'b001110100111;
		16'b1100101001111110: color_data = 12'b001110100111;
		16'b1100101001111111: color_data = 12'b001110100111;
		16'b1100101010000000: color_data = 12'b001110100111;
		16'b1100101010001101: color_data = 12'b001110100111;
		16'b1100101010001110: color_data = 12'b001110100111;
		16'b1100101010001111: color_data = 12'b001110100111;
		16'b1100101010010000: color_data = 12'b001110100111;
		16'b1100101010010001: color_data = 12'b001110100111;
		16'b1100101010010010: color_data = 12'b001110100111;
		16'b1100101010010011: color_data = 12'b001110100111;
		16'b1100101010010100: color_data = 12'b001110100111;
		16'b1100101010010101: color_data = 12'b001110100111;
		16'b1100101010010110: color_data = 12'b001110100111;
		16'b1100101010010111: color_data = 12'b001110100111;
		16'b1100101010011000: color_data = 12'b001110100111;
		16'b1100101010011001: color_data = 12'b001110100111;
		16'b1100101010100000: color_data = 12'b001110100111;
		16'b1100101010100001: color_data = 12'b001110100111;
		16'b1100101010100010: color_data = 12'b001110100111;
		16'b1100101010100011: color_data = 12'b001110100111;
		16'b1100101010100100: color_data = 12'b001110100111;
		16'b1100101010100101: color_data = 12'b001110100111;
		16'b1100101010100110: color_data = 12'b001110100111;
		16'b1100101010100111: color_data = 12'b001110100111;
		16'b1100101010101000: color_data = 12'b001110100111;
		16'b1100101010101001: color_data = 12'b001110100111;
		16'b1100101010101010: color_data = 12'b001110100111;
		16'b1100101010101011: color_data = 12'b001110100111;
		16'b1100101010101100: color_data = 12'b001110100111;
		16'b1100101010101101: color_data = 12'b001110100111;
		16'b1100101010101110: color_data = 12'b001110100111;
		16'b1100101010101111: color_data = 12'b001110100111;
		16'b1100101010110000: color_data = 12'b001110100111;
		16'b1100101010110001: color_data = 12'b001110100111;
		16'b1100101010110010: color_data = 12'b001110100111;
		16'b1100101010110011: color_data = 12'b001110100111;
		16'b1100101010110100: color_data = 12'b001110100111;
		16'b1100101010110101: color_data = 12'b001110100111;
		16'b1100101010110110: color_data = 12'b001110100111;
		16'b1100101010110111: color_data = 12'b001110100111;
		16'b1100101010111000: color_data = 12'b001110100111;
		16'b1100101010111001: color_data = 12'b001110100111;
		16'b1100101010111010: color_data = 12'b001110100111;
		16'b1100101010111011: color_data = 12'b001110100111;
		16'b1100101010111100: color_data = 12'b001110100111;
		16'b1100101010111101: color_data = 12'b001110100111;
		16'b1100101010111110: color_data = 12'b001110100111;
		16'b1100101010111111: color_data = 12'b001110100111;
		16'b1100101011000000: color_data = 12'b001110100111;
		16'b1100101011000001: color_data = 12'b001110100111;
		16'b1100101011000010: color_data = 12'b001110100111;
		16'b1100101011000011: color_data = 12'b001110100111;
		16'b1100101011000100: color_data = 12'b001110100111;
		16'b1100101011001011: color_data = 12'b001110100111;
		16'b1100101011001100: color_data = 12'b001110100111;
		16'b1100101011001101: color_data = 12'b001110100111;
		16'b1100101011001110: color_data = 12'b001110100111;
		16'b1100101011001111: color_data = 12'b001110100111;
		16'b1100101011010000: color_data = 12'b001110100111;
		16'b1100101011010001: color_data = 12'b001110100111;
		16'b1100101011010010: color_data = 12'b001110100111;
		16'b1100101011010011: color_data = 12'b001110100111;
		16'b1100101011010100: color_data = 12'b001110100111;
		16'b1100101011010101: color_data = 12'b001110100111;
		16'b1100101011010110: color_data = 12'b001110100111;
		16'b1100101011111100: color_data = 12'b001110100111;
		16'b1100101011111101: color_data = 12'b001110100111;
		16'b1100101011111110: color_data = 12'b001110100111;
		16'b1100101011111111: color_data = 12'b001110100111;
		16'b1100101100000000: color_data = 12'b001110100111;
		16'b1100101100000001: color_data = 12'b001110100111;
		16'b1100101100000010: color_data = 12'b001110100111;
		16'b1100101100000011: color_data = 12'b001110100111;
		16'b1100101100000100: color_data = 12'b001110100111;
		16'b1100101100000101: color_data = 12'b001110100111;
		16'b1100101100000110: color_data = 12'b001110100111;
		16'b1100101100000111: color_data = 12'b001110100111;
		16'b1100101100001000: color_data = 12'b001110100111;
		16'b1100101100001001: color_data = 12'b001110100111;
		16'b1100101100001010: color_data = 12'b001110100111;
		16'b1100101100001011: color_data = 12'b001110100111;
		16'b1100101100001100: color_data = 12'b001110100111;
		16'b1100101100001101: color_data = 12'b001110100111;
		16'b1100101100001110: color_data = 12'b001110100111;
		16'b1100101100001111: color_data = 12'b001110100111;
		16'b1100101100010000: color_data = 12'b001110100111;
		16'b1100101100010001: color_data = 12'b001110100111;
		16'b1100101100010010: color_data = 12'b001110100111;
		16'b1100101100010011: color_data = 12'b001110100111;
		16'b1100101100010100: color_data = 12'b001110100111;
		16'b1100101100010101: color_data = 12'b001110100111;
		16'b1100101100010110: color_data = 12'b001110100111;
		16'b1100101100010111: color_data = 12'b001110100111;
		16'b1100101100011000: color_data = 12'b001110100111;
		16'b1100101100011001: color_data = 12'b001110100111;
		16'b1100101100011010: color_data = 12'b001110100111;
		16'b1100101100011011: color_data = 12'b001110100111;
		16'b1100101100011100: color_data = 12'b001110100111;
		16'b1100101100011101: color_data = 12'b001110100111;
		16'b1100101100011110: color_data = 12'b001110100111;
		16'b1100101100011111: color_data = 12'b001110100111;
		16'b1100101100100000: color_data = 12'b001110100111;
		16'b1100101100101101: color_data = 12'b001110100111;
		16'b1100101100101110: color_data = 12'b001110100111;
		16'b1100101100101111: color_data = 12'b001110100111;
		16'b1100101100110000: color_data = 12'b001110100111;
		16'b1100101100110001: color_data = 12'b001110100111;
		16'b1100101100110010: color_data = 12'b001110100111;
		16'b1100101100110011: color_data = 12'b001110100111;
		16'b1100101100110100: color_data = 12'b001110100111;
		16'b1100101100110101: color_data = 12'b001110100111;
		16'b1100101100110110: color_data = 12'b001110100111;
		16'b1100101100110111: color_data = 12'b001110100111;
		16'b1100101100111000: color_data = 12'b001110100111;
		16'b1100101101000101: color_data = 12'b001110100111;
		16'b1100101101000110: color_data = 12'b001110100111;
		16'b1100101101000111: color_data = 12'b001110100111;
		16'b1100101101001000: color_data = 12'b001110100111;
		16'b1100101101001001: color_data = 12'b001110100111;
		16'b1100101101001010: color_data = 12'b001110100111;
		16'b1100101101001011: color_data = 12'b001110100111;
		16'b1100101101001100: color_data = 12'b001110100111;
		16'b1100101101001101: color_data = 12'b001110100111;
		16'b1100101101001110: color_data = 12'b001110100111;
		16'b1100101101001111: color_data = 12'b001110100111;
		16'b1100101101010000: color_data = 12'b001110100111;
		16'b1100101101010001: color_data = 12'b001110100111;
		16'b1100101101011000: color_data = 12'b001110100111;
		16'b1100101101011001: color_data = 12'b001110100111;
		16'b1100101101011010: color_data = 12'b001110100111;
		16'b1100101101011011: color_data = 12'b001110100111;
		16'b1100101101011100: color_data = 12'b001110100111;
		16'b1100101101011101: color_data = 12'b001110100111;
		16'b1100101101011110: color_data = 12'b001110100111;
		16'b1100101101011111: color_data = 12'b001110100111;
		16'b1100101101100000: color_data = 12'b001110100111;
		16'b1100101101100001: color_data = 12'b001110100111;
		16'b1100101101100010: color_data = 12'b001110100111;
		16'b1100101101100011: color_data = 12'b001110100111;
		16'b1100101101100100: color_data = 12'b001110100111;
		16'b1100101101100101: color_data = 12'b001110100111;
		16'b1100101101100110: color_data = 12'b001110100111;
		16'b1100101101100111: color_data = 12'b001110100111;
		16'b1100101101101000: color_data = 12'b001110100111;
		16'b1100101101101001: color_data = 12'b001110100111;
		16'b1100101101101010: color_data = 12'b001110100111;
		16'b1100101101101011: color_data = 12'b001110100111;
		16'b1100101101101100: color_data = 12'b001110100111;
		16'b1100101101101101: color_data = 12'b001110100111;
		16'b1100101101101110: color_data = 12'b001110100111;
		16'b1100101101101111: color_data = 12'b001110100111;
		16'b1100101101110000: color_data = 12'b001110100111;
		16'b1100101101110001: color_data = 12'b001110100111;
		16'b1100101101110010: color_data = 12'b001110100111;
		16'b1100101101110011: color_data = 12'b001110100111;
		16'b1100101101110100: color_data = 12'b001110100111;
		16'b1100101101110101: color_data = 12'b001110100111;
		16'b1100101101110110: color_data = 12'b001110100111;
		16'b1100101101110111: color_data = 12'b001110100111;
		16'b1100101101111000: color_data = 12'b001110100111;
		16'b1100101101111001: color_data = 12'b001110100111;
		16'b1100101101111010: color_data = 12'b001110100111;
		16'b1100101101111011: color_data = 12'b001110100111;


    default: color_data = 12'b000000000000;
	endcase
endmodule