module no_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		11'b00000000000: color_data = 12'b110011110111;
		11'b00000000001: color_data = 12'b110011110111;
		11'b00000000010: color_data = 12'b110011110111;
		11'b00000000011: color_data = 12'b110011110111;
		11'b00000001101: color_data = 12'b110011110111;
		11'b00000001110: color_data = 12'b110011110111;
		11'b00000001111: color_data = 12'b110011110111;
		11'b00000010000: color_data = 12'b110011110111;
		11'b00000010001: color_data = 12'b110011110111;
		11'b00000010101: color_data = 12'b110011110111;
		11'b00000010110: color_data = 12'b110011110111;
		11'b00000010111: color_data = 12'b110011110111;
		11'b00000011000: color_data = 12'b110011110111;
		11'b00000011001: color_data = 12'b110011110111;
		11'b00000011010: color_data = 12'b110011110111;
		11'b00000011011: color_data = 12'b110011110111;
		11'b00000011100: color_data = 12'b110011110111;
		11'b00000011101: color_data = 12'b110011110111;
		11'b00000011110: color_data = 12'b110011110111;
		11'b00000011111: color_data = 12'b110011110111;
		11'b00001000000: color_data = 12'b110011110111;
		11'b00001000001: color_data = 12'b110011110111;
		11'b00001000010: color_data = 12'b110011110111;
		11'b00001000011: color_data = 12'b110011110111;
		11'b00001001101: color_data = 12'b110011110111;
		11'b00001001110: color_data = 12'b110011110111;
		11'b00001010001: color_data = 12'b110011110111;
		11'b00001010100: color_data = 12'b110011110111;
		11'b00001010101: color_data = 12'b110011110111;
		11'b00001010110: color_data = 12'b110011110111;
		11'b00001011101: color_data = 12'b110011110111;
		11'b00001011110: color_data = 12'b110011110111;
		11'b00001011111: color_data = 12'b110011110111;
		11'b00001100000: color_data = 12'b110011110111;
		11'b00010000000: color_data = 12'b110011110111;
		11'b00010000001: color_data = 12'b110011110111;
		11'b00010000010: color_data = 12'b110011110111;
		11'b00010000011: color_data = 12'b110011110111;
		11'b00010000100: color_data = 12'b110011110111;
		11'b00010001101: color_data = 12'b110011110111;
		11'b00010001110: color_data = 12'b110011110111;
		11'b00010010001: color_data = 12'b110011110111;
		11'b00010010011: color_data = 12'b110011110111;
		11'b00010010100: color_data = 12'b110011110111;
		11'b00010010101: color_data = 12'b110011110111;
		11'b00010011101: color_data = 12'b110011110111;
		11'b00010011111: color_data = 12'b110011110111;
		11'b00010100000: color_data = 12'b110011110111;
		11'b00010100001: color_data = 12'b110011110111;
		11'b00011000000: color_data = 12'b110011110111;
		11'b00011000001: color_data = 12'b110011110111;
		11'b00011000011: color_data = 12'b110011110111;
		11'b00011000100: color_data = 12'b110011110111;
		11'b00011000101: color_data = 12'b110011110111;
		11'b00011001101: color_data = 12'b110011110111;
		11'b00011001110: color_data = 12'b110011110111;
		11'b00011010001: color_data = 12'b110011110111;
		11'b00011010011: color_data = 12'b110011110111;
		11'b00011010100: color_data = 12'b110011110111;
		11'b00011010101: color_data = 12'b110011110111;
		11'b00011011101: color_data = 12'b110011110111;
		11'b00011011111: color_data = 12'b110011110111;
		11'b00011100000: color_data = 12'b110011110111;
		11'b00011100001: color_data = 12'b110011110111;
		11'b00100000000: color_data = 12'b110011110111;
		11'b00100000001: color_data = 12'b110011110111;
		11'b00100000011: color_data = 12'b110011110111;
		11'b00100000100: color_data = 12'b110011110111;
		11'b00100000101: color_data = 12'b110011110111;
		11'b00100001101: color_data = 12'b110011110111;
		11'b00100001110: color_data = 12'b110011110111;
		11'b00100010001: color_data = 12'b110011110111;
		11'b00100010011: color_data = 12'b110011110111;
		11'b00100010100: color_data = 12'b110011110111;
		11'b00100010101: color_data = 12'b110011110111;
		11'b00100011101: color_data = 12'b110011110111;
		11'b00100011111: color_data = 12'b110011110111;
		11'b00100100000: color_data = 12'b110011110111;
		11'b00100100001: color_data = 12'b110011110111;
		11'b00101000000: color_data = 12'b110011110111;
		11'b00101000001: color_data = 12'b110011110111;
		11'b00101000011: color_data = 12'b110011110111;
		11'b00101000100: color_data = 12'b110011110111;
		11'b00101000101: color_data = 12'b110011110111;
		11'b00101000110: color_data = 12'b110011110111;
		11'b00101001101: color_data = 12'b110011110111;
		11'b00101001110: color_data = 12'b110011110111;
		11'b00101010001: color_data = 12'b110011110111;
		11'b00101010011: color_data = 12'b110011110111;
		11'b00101010100: color_data = 12'b110011110111;
		11'b00101010101: color_data = 12'b110011110111;
		11'b00101011101: color_data = 12'b110011110111;
		11'b00101011111: color_data = 12'b110011110111;
		11'b00101100000: color_data = 12'b110011110111;
		11'b00101100001: color_data = 12'b110011110111;
		11'b00110000000: color_data = 12'b110011110111;
		11'b00110000001: color_data = 12'b110011110111;
		11'b00110000011: color_data = 12'b110011110111;
		11'b00110000100: color_data = 12'b110011110111;
		11'b00110000101: color_data = 12'b110011110111;
		11'b00110000110: color_data = 12'b110011110111;
		11'b00110001101: color_data = 12'b110011110111;
		11'b00110001110: color_data = 12'b110011110111;
		11'b00110010001: color_data = 12'b110011110111;
		11'b00110010011: color_data = 12'b110011110111;
		11'b00110010100: color_data = 12'b110011110111;
		11'b00110010101: color_data = 12'b110011110111;
		11'b00110011101: color_data = 12'b110011110111;
		11'b00110011111: color_data = 12'b110011110111;
		11'b00110100000: color_data = 12'b110011110111;
		11'b00110100001: color_data = 12'b110011110111;
		11'b00111000000: color_data = 12'b110011110111;
		11'b00111000001: color_data = 12'b110011110111;
		11'b00111000011: color_data = 12'b110011110111;
		11'b00111000101: color_data = 12'b110011110111;
		11'b00111000110: color_data = 12'b110011110111;
		11'b00111000111: color_data = 12'b110011110111;
		11'b00111001101: color_data = 12'b110011110111;
		11'b00111001110: color_data = 12'b110011110111;
		11'b00111010001: color_data = 12'b110011110111;
		11'b00111010011: color_data = 12'b110011110111;
		11'b00111010100: color_data = 12'b110011110111;
		11'b00111010101: color_data = 12'b110011110111;
		11'b00111011101: color_data = 12'b110011110111;
		11'b00111011111: color_data = 12'b110011110111;
		11'b00111100000: color_data = 12'b110011110111;
		11'b00111100001: color_data = 12'b110011110111;
		11'b01000000000: color_data = 12'b110011110111;
		11'b01000000001: color_data = 12'b110011110111;
		11'b01000000011: color_data = 12'b110011110111;
		11'b01000000110: color_data = 12'b110011110111;
		11'b01000000111: color_data = 12'b110011110111;
		11'b01000001000: color_data = 12'b110011110111;
		11'b01000001101: color_data = 12'b110011110111;
		11'b01000001110: color_data = 12'b110011110111;
		11'b01000010001: color_data = 12'b110011110111;
		11'b01000010011: color_data = 12'b110011110111;
		11'b01000010100: color_data = 12'b110011110111;
		11'b01000010101: color_data = 12'b110011110111;
		11'b01000011101: color_data = 12'b110011110111;
		11'b01000011111: color_data = 12'b110011110111;
		11'b01000100000: color_data = 12'b110011110111;
		11'b01000100001: color_data = 12'b110011110111;
		11'b01001000000: color_data = 12'b110011110111;
		11'b01001000001: color_data = 12'b110011110111;
		11'b01001000011: color_data = 12'b110011110111;
		11'b01001000110: color_data = 12'b110011110111;
		11'b01001000111: color_data = 12'b110011110111;
		11'b01001001000: color_data = 12'b110011110111;
		11'b01001001101: color_data = 12'b110011110111;
		11'b01001001110: color_data = 12'b110011110111;
		11'b01001010001: color_data = 12'b110011110111;
		11'b01001010011: color_data = 12'b110011110111;
		11'b01001010100: color_data = 12'b110011110111;
		11'b01001010101: color_data = 12'b110011110111;
		11'b01001011101: color_data = 12'b110011110111;
		11'b01001011111: color_data = 12'b110011110111;
		11'b01001100000: color_data = 12'b110011110111;
		11'b01001100001: color_data = 12'b110011110111;
		11'b01010000000: color_data = 12'b110011110111;
		11'b01010000001: color_data = 12'b110011110111;
		11'b01010000011: color_data = 12'b110011110111;
		11'b01010000111: color_data = 12'b110011110111;
		11'b01010001000: color_data = 12'b110011110111;
		11'b01010001001: color_data = 12'b110011110111;
		11'b01010001101: color_data = 12'b110011110111;
		11'b01010001110: color_data = 12'b110011110111;
		11'b01010010001: color_data = 12'b110011110111;
		11'b01010010011: color_data = 12'b110011110111;
		11'b01010010100: color_data = 12'b110011110111;
		11'b01010010101: color_data = 12'b110011110111;
		11'b01010011101: color_data = 12'b110011110111;
		11'b01010011111: color_data = 12'b110011110111;
		11'b01010100000: color_data = 12'b110011110111;
		11'b01010100001: color_data = 12'b110011110111;
		11'b01011000000: color_data = 12'b110011110111;
		11'b01011000001: color_data = 12'b110011110111;
		11'b01011000011: color_data = 12'b110011110111;
		11'b01011001000: color_data = 12'b110011110111;
		11'b01011001001: color_data = 12'b110011110111;
		11'b01011001010: color_data = 12'b110011110111;
		11'b01011001101: color_data = 12'b110011110111;
		11'b01011001110: color_data = 12'b110011110111;
		11'b01011010001: color_data = 12'b110011110111;
		11'b01011010011: color_data = 12'b110011110111;
		11'b01011010100: color_data = 12'b110011110111;
		11'b01011010101: color_data = 12'b110011110111;
		11'b01011011101: color_data = 12'b110011110111;
		11'b01011011111: color_data = 12'b110011110111;
		11'b01011100000: color_data = 12'b110011110111;
		11'b01011100001: color_data = 12'b110011110111;
		11'b01100000000: color_data = 12'b110011110111;
		11'b01100000001: color_data = 12'b110011110111;
		11'b01100000011: color_data = 12'b110011110111;
		11'b01100001000: color_data = 12'b110011110111;
		11'b01100001001: color_data = 12'b110011110111;
		11'b01100001010: color_data = 12'b110011110111;
		11'b01100001101: color_data = 12'b110011110111;
		11'b01100001110: color_data = 12'b110011110111;
		11'b01100010001: color_data = 12'b110011110111;
		11'b01100010011: color_data = 12'b110011110111;
		11'b01100010100: color_data = 12'b110011110111;
		11'b01100010101: color_data = 12'b110011110111;
		11'b01100011101: color_data = 12'b110011110111;
		11'b01100011111: color_data = 12'b110011110111;
		11'b01100100000: color_data = 12'b110011110111;
		11'b01100100001: color_data = 12'b110011110111;
		11'b01101000000: color_data = 12'b110011110111;
		11'b01101000001: color_data = 12'b110011110111;
		11'b01101000011: color_data = 12'b110011110111;
		11'b01101001001: color_data = 12'b110011110111;
		11'b01101001010: color_data = 12'b110011110111;
		11'b01101001011: color_data = 12'b110011110111;
		11'b01101001101: color_data = 12'b110011110111;
		11'b01101001110: color_data = 12'b110011110111;
		11'b01101010001: color_data = 12'b110011110111;
		11'b01101010011: color_data = 12'b110011110111;
		11'b01101010100: color_data = 12'b110011110111;
		11'b01101010101: color_data = 12'b110011110111;
		11'b01101011101: color_data = 12'b110011110111;
		11'b01101011111: color_data = 12'b110011110111;
		11'b01101100000: color_data = 12'b110011110111;
		11'b01101100001: color_data = 12'b110011110111;
		11'b01110000000: color_data = 12'b110011110111;
		11'b01110000001: color_data = 12'b110011110111;
		11'b01110000011: color_data = 12'b110011110111;
		11'b01110001010: color_data = 12'b110011110111;
		11'b01110001011: color_data = 12'b110011110111;
		11'b01110001100: color_data = 12'b110011110111;
		11'b01110001101: color_data = 12'b110011110111;
		11'b01110001110: color_data = 12'b110011110111;
		11'b01110010001: color_data = 12'b110011110111;
		11'b01110010011: color_data = 12'b110011110111;
		11'b01110010100: color_data = 12'b110011110111;
		11'b01110010101: color_data = 12'b110011110111;
		11'b01110011101: color_data = 12'b110011110111;
		11'b01110011111: color_data = 12'b110011110111;
		11'b01110100000: color_data = 12'b110011110111;
		11'b01110100001: color_data = 12'b110011110111;
		11'b01111000000: color_data = 12'b110011110111;
		11'b01111000001: color_data = 12'b110011110111;
		11'b01111000011: color_data = 12'b110011110111;
		11'b01111001010: color_data = 12'b110011110111;
		11'b01111001011: color_data = 12'b110011110111;
		11'b01111001100: color_data = 12'b110011110111;
		11'b01111001101: color_data = 12'b110011110111;
		11'b01111001110: color_data = 12'b110011110111;
		11'b01111010001: color_data = 12'b110011110111;
		11'b01111010100: color_data = 12'b110011110111;
		11'b01111010101: color_data = 12'b110011110111;
		11'b01111010110: color_data = 12'b110011110111;
		11'b01111011101: color_data = 12'b110011110111;
		11'b01111011110: color_data = 12'b110011110111;
		11'b01111011111: color_data = 12'b110011110111;
		11'b01111100000: color_data = 12'b110011110111;
		11'b10000000000: color_data = 12'b110011110111;
		11'b10000000001: color_data = 12'b110011110111;
		11'b10000000010: color_data = 12'b110011110111;
		11'b10000000011: color_data = 12'b110011110111;
		11'b10000001011: color_data = 12'b110011110111;
		11'b10000001100: color_data = 12'b110011110111;
		11'b10000001101: color_data = 12'b110011110111;
		11'b10000001110: color_data = 12'b110011110111;
		11'b10000001111: color_data = 12'b110011110111;
		11'b10000010000: color_data = 12'b110011110111;
		11'b10000010001: color_data = 12'b110011110111;
		11'b10000010101: color_data = 12'b110011110111;
		11'b10000010110: color_data = 12'b110011110111;
		11'b10000010111: color_data = 12'b110011110111;
		11'b10000011000: color_data = 12'b110011110111;
		11'b10000011001: color_data = 12'b110011110111;
		11'b10000011010: color_data = 12'b110011110111;
		11'b10000011011: color_data = 12'b110011110111;
		11'b10000011100: color_data = 12'b110011110111;
		11'b10000011101: color_data = 12'b110011110111;
		11'b10000011110: color_data = 12'b110011110111;
		11'b10000011111: color_data = 12'b110011110111;
		11'b10001000000: color_data = 12'b110011110111;
		11'b10001000001: color_data = 12'b110011110111;
		11'b10001000010: color_data = 12'b110011110111;
		11'b10001000011: color_data = 12'b110011110111;
		11'b10001001011: color_data = 12'b110011110111;
		11'b10001001100: color_data = 12'b110011110111;
		11'b10001001101: color_data = 12'b110011110111;
		11'b10001001110: color_data = 12'b110011110111;
		11'b10001001111: color_data = 12'b110011110111;
		11'b10001010000: color_data = 12'b110011110111;
		11'b10001010001: color_data = 12'b110011110111;
		11'b10001010110: color_data = 12'b110011110111;
		11'b10001010111: color_data = 12'b110011110111;
		11'b10001011000: color_data = 12'b110011110111;
		11'b10001011001: color_data = 12'b110011110111;
		11'b10001011010: color_data = 12'b110011110111;
		11'b10001011011: color_data = 12'b110011110111;
		11'b10001011100: color_data = 12'b110011110111;
		11'b10001011101: color_data = 12'b110011110111;
		11'b10001011110: color_data = 12'b110011110111;
        default: color_data = 12'b000000000000;
	endcase
endmodule