module heart_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
				10'b0000000100: color_data = 12'b011011111110;
		10'b0000000101: color_data = 12'b011011111110;
		10'b0000000110: color_data = 12'b011011111110;
		10'b0000000111: color_data = 12'b011011111110;
		10'b0000001000: color_data = 12'b011011111110;
		10'b0000001001: color_data = 12'b011011111110;
		10'b0000010000: color_data = 12'b011011111110;
		10'b0000010001: color_data = 12'b011011111110;
		10'b0000010010: color_data = 12'b011011111110;
		10'b0000010011: color_data = 12'b011011111110;
		10'b0000010100: color_data = 12'b011011111110;
		10'b0000010101: color_data = 12'b011011111110;
		10'b0000100010: color_data = 12'b011011111110;
		10'b0000100011: color_data = 12'b011011111110;
		10'b0000100100: color_data = 12'b101100010010;
		10'b0000100101: color_data = 12'b101100010010;
		10'b0000100110: color_data = 12'b101100010010;
		10'b0000100111: color_data = 12'b101100010010;
		10'b0000101000: color_data = 12'b101100010010;
		10'b0000101001: color_data = 12'b101100010010;
		10'b0000101010: color_data = 12'b011011111110;
		10'b0000101011: color_data = 12'b011011111110;
		10'b0000101110: color_data = 12'b011011111110;
		10'b0000101111: color_data = 12'b011011111110;
		10'b0000110000: color_data = 12'b101100010011;
		10'b0000110001: color_data = 12'b110000010010;
		10'b0000110010: color_data = 12'b101100010010;
		10'b0000110011: color_data = 12'b101100010010;
		10'b0000110100: color_data = 12'b101100010010;
		10'b0000110101: color_data = 12'b101100010010;
		10'b0000110110: color_data = 12'b011011111110;
		10'b0000110111: color_data = 12'b011011111110;
		10'b0001000010: color_data = 12'b011011111110;
		10'b0001000011: color_data = 12'b011011111110;
		10'b0001000100: color_data = 12'b101100010010;
		10'b0001000101: color_data = 12'b101100010010;
		10'b0001000110: color_data = 12'b101100010010;
		10'b0001000111: color_data = 12'b101100010010;
		10'b0001001000: color_data = 12'b101100010010;
		10'b0001001001: color_data = 12'b101100010011;
		10'b0001001010: color_data = 12'b011011111110;
		10'b0001001011: color_data = 12'b011011111110;
		10'b0001001110: color_data = 12'b011011111110;
		10'b0001001111: color_data = 12'b011011111110;
		10'b0001010000: color_data = 12'b101100010011;
		10'b0001010001: color_data = 12'b101100010010;
		10'b0001010010: color_data = 12'b101100010010;
		10'b0001010011: color_data = 12'b101100010010;
		10'b0001010100: color_data = 12'b101100010010;
		10'b0001010101: color_data = 12'b101100100010;
		10'b0001010110: color_data = 12'b011011111110;
		10'b0001010111: color_data = 12'b011011111110;
		10'b0001100001: color_data = 12'b000100000000;
		10'b0001100010: color_data = 12'b011011111110;
		10'b0001100011: color_data = 12'b011011111110;
		10'b0001100100: color_data = 12'b101100010011;
		10'b0001100101: color_data = 12'b101100010010;
		10'b0001100110: color_data = 12'b101100010010;
		10'b0001100111: color_data = 12'b101100100011;
		10'b0001101000: color_data = 12'b101100010010;
		10'b0001101001: color_data = 12'b101100100010;
		10'b0001101010: color_data = 12'b011011111110;
		10'b0001101011: color_data = 12'b011011111110;
		10'b0001101110: color_data = 12'b011011111110;
		10'b0001101111: color_data = 12'b011011111110;
		10'b0001110000: color_data = 12'b110000010011;
		10'b0001110001: color_data = 12'b110000010010;
		10'b0001110010: color_data = 12'b101100010010;
		10'b0001110011: color_data = 12'b101100010010;
		10'b0001110100: color_data = 12'b101100010010;
		10'b0001110101: color_data = 12'b101100100011;
		10'b0001110110: color_data = 12'b011011111110;
		10'b0001110111: color_data = 12'b011011111110;
		10'b0010000000: color_data = 12'b011011111110;
		10'b0010000001: color_data = 12'b011011111110;
		10'b0010000010: color_data = 12'b110000010011;
		10'b0010000011: color_data = 12'b110000010011;
		10'b0010000100: color_data = 12'b111111111111;
		10'b0010000101: color_data = 12'b111111111111;
		10'b0010000110: color_data = 12'b111111111111;
		10'b0010000111: color_data = 12'b111111111111;
		10'b0010001000: color_data = 12'b110000010010;
		10'b0010001001: color_data = 12'b110000010011;
		10'b0010001010: color_data = 12'b110000010010;
		10'b0010001011: color_data = 12'b101100010010;
		10'b0010001100: color_data = 12'b011011111110;
		10'b0010001101: color_data = 12'b011011111110;
		10'b0010001110: color_data = 12'b101100100011;
		10'b0010001111: color_data = 12'b110000010010;
		10'b0010010000: color_data = 12'b110000010010;
		10'b0010010001: color_data = 12'b101100010010;
		10'b0010010010: color_data = 12'b101100010010;
		10'b0010010011: color_data = 12'b101100010010;
		10'b0010010100: color_data = 12'b101100010010;
		10'b0010010101: color_data = 12'b110000010010;
		10'b0010010110: color_data = 12'b110000010010;
		10'b0010010111: color_data = 12'b101100100010;
		10'b0010011000: color_data = 12'b011011111110;
		10'b0010011001: color_data = 12'b011011111110;
		10'b0010100000: color_data = 12'b011011111110;
		10'b0010100001: color_data = 12'b011011111110;
		10'b0010100010: color_data = 12'b101100010010;
		10'b0010100011: color_data = 12'b110000010010;
		10'b0010100100: color_data = 12'b111111111111;
		10'b0010100101: color_data = 12'b011011111110;
		10'b0010100110: color_data = 12'b011011111110;
		10'b0010100111: color_data = 12'b111111111111;
		10'b0010101000: color_data = 12'b110000010010;
		10'b0010101001: color_data = 12'b101100100011;
		10'b0010101010: color_data = 12'b101100100011;
		10'b0010101011: color_data = 12'b101100100011;
		10'b0010101100: color_data = 12'b011011111110;
		10'b0010101101: color_data = 12'b011011111110;
		10'b0010101110: color_data = 12'b101100010011;
		10'b0010101111: color_data = 12'b110000010011;
		10'b0010110000: color_data = 12'b110000010011;
		10'b0010110001: color_data = 12'b110000010010;
		10'b0010110010: color_data = 12'b101100010010;
		10'b0010110011: color_data = 12'b101100010010;
		10'b0010110100: color_data = 12'b101100010010;
		10'b0010110101: color_data = 12'b101100010010;
		10'b0010110110: color_data = 12'b101100010010;
		10'b0010110111: color_data = 12'b101100010011;
		10'b0010111000: color_data = 12'b011011111110;
		10'b0010111001: color_data = 12'b011011111110;
		10'b0011000000: color_data = 12'b011011111110;
		10'b0011000001: color_data = 12'b011011111110;
		10'b0011000010: color_data = 12'b101100010010;
		10'b0011000011: color_data = 12'b101100010011;
		10'b0011000100: color_data = 12'b111111111111;
		10'b0011000101: color_data = 12'b111111001100;
		10'b0011000110: color_data = 12'b101100010011;
		10'b0011000111: color_data = 12'b101100010011;
		10'b0011001000: color_data = 12'b110000100010;
		10'b0011001001: color_data = 12'b101100010010;
		10'b0011001010: color_data = 12'b101100100010;
		10'b0011001011: color_data = 12'b110000010010;
		10'b0011001100: color_data = 12'b101100100010;
		10'b0011001101: color_data = 12'b101100100011;
		10'b0011001110: color_data = 12'b101100010010;
		10'b0011001111: color_data = 12'b101100010010;
		10'b0011010000: color_data = 12'b101100010010;
		10'b0011010001: color_data = 12'b101100010010;
		10'b0011010010: color_data = 12'b101100010010;
		10'b0011010011: color_data = 12'b101100010010;
		10'b0011010100: color_data = 12'b101100010010;
		10'b0011010101: color_data = 12'b101100010010;
		10'b0011010110: color_data = 12'b101100010010;
		10'b0011010111: color_data = 12'b110000010010;
		10'b0011011000: color_data = 12'b011011111110;
		10'b0011011001: color_data = 12'b011011111110;
		10'b0011100000: color_data = 12'b011011111110;
		10'b0011100001: color_data = 12'b011011111110;
		10'b0011100010: color_data = 12'b101100010010;
		10'b0011100011: color_data = 12'b101100010011;
		10'b0011100100: color_data = 12'b111111111111;
		10'b0011100101: color_data = 12'b111111001101;
		10'b0011100110: color_data = 12'b110000010010;
		10'b0011100111: color_data = 12'b101100010010;
		10'b0011101000: color_data = 12'b101100010010;
		10'b0011101001: color_data = 12'b101100010010;
		10'b0011101010: color_data = 12'b101100010010;
		10'b0011101011: color_data = 12'b101100010010;
		10'b0011101100: color_data = 12'b101100010010;
		10'b0011101101: color_data = 12'b101100010010;
		10'b0011101110: color_data = 12'b101100010010;
		10'b0011101111: color_data = 12'b101100010010;
		10'b0011110000: color_data = 12'b101100010010;
		10'b0011110001: color_data = 12'b101100010010;
		10'b0011110010: color_data = 12'b101100010010;
		10'b0011110011: color_data = 12'b101100010010;
		10'b0011110100: color_data = 12'b101100010010;
		10'b0011110101: color_data = 12'b101100010010;
		10'b0011110110: color_data = 12'b101100010010;
		10'b0011110111: color_data = 12'b110000010010;
		10'b0011111000: color_data = 12'b011011111110;
		10'b0011111001: color_data = 12'b011011111110;
		10'b0100000000: color_data = 12'b011011111110;
		10'b0100000001: color_data = 12'b011011111110;
		10'b0100000010: color_data = 12'b101100010010;
		10'b0100000011: color_data = 12'b101100010011;
		10'b0100000100: color_data = 12'b101100010010;
		10'b0100000101: color_data = 12'b110000010010;
		10'b0100000110: color_data = 12'b101100010011;
		10'b0100000111: color_data = 12'b101100010010;
		10'b0100001000: color_data = 12'b101100010010;
		10'b0100001001: color_data = 12'b101100010010;
		10'b0100001010: color_data = 12'b101100010010;
		10'b0100001011: color_data = 12'b101100010010;
		10'b0100001100: color_data = 12'b101100010010;
		10'b0100001101: color_data = 12'b101100010010;
		10'b0100001110: color_data = 12'b101100010010;
		10'b0100001111: color_data = 12'b101100010010;
		10'b0100010000: color_data = 12'b101100010010;
		10'b0100010001: color_data = 12'b101100010010;
		10'b0100010010: color_data = 12'b101100010010;
		10'b0100010011: color_data = 12'b101100010010;
		10'b0100010100: color_data = 12'b101100010010;
		10'b0100010101: color_data = 12'b101100010010;
		10'b0100010110: color_data = 12'b101100010010;
		10'b0100010111: color_data = 12'b110000010010;
		10'b0100011000: color_data = 12'b011011111110;
		10'b0100011001: color_data = 12'b011011111110;
		10'b0100100000: color_data = 12'b011011111110;
		10'b0100100001: color_data = 12'b011011111110;
		10'b0100100010: color_data = 12'b101100010011;
		10'b0100100011: color_data = 12'b110000010011;
		10'b0100100100: color_data = 12'b101100010011;
		10'b0100100101: color_data = 12'b101100010010;
		10'b0100100110: color_data = 12'b101100010010;
		10'b0100100111: color_data = 12'b101100010010;
		10'b0100101000: color_data = 12'b101100010010;
		10'b0100101001: color_data = 12'b101100010010;
		10'b0100101010: color_data = 12'b101100010010;
		10'b0100101011: color_data = 12'b101100010010;
		10'b0100101100: color_data = 12'b101100010010;
		10'b0100101101: color_data = 12'b101100010010;
		10'b0100101110: color_data = 12'b101100010010;
		10'b0100101111: color_data = 12'b101100010010;
		10'b0100110000: color_data = 12'b101100010010;
		10'b0100110001: color_data = 12'b101100010010;
		10'b0100110010: color_data = 12'b101100010010;
		10'b0100110011: color_data = 12'b101100010010;
		10'b0100110100: color_data = 12'b101100010010;
		10'b0100110101: color_data = 12'b101100100010;
		10'b0100110110: color_data = 12'b110000010010;
		10'b0100110111: color_data = 12'b101100010011;
		10'b0100111000: color_data = 12'b011011111110;
		10'b0100111001: color_data = 12'b011011111110;
		10'b0101000010: color_data = 12'b011011111110;
		10'b0101000011: color_data = 12'b011011111110;
		10'b0101000100: color_data = 12'b101100100010;
		10'b0101000101: color_data = 12'b101100010010;
		10'b0101000110: color_data = 12'b101100010010;
		10'b0101000111: color_data = 12'b101100010010;
		10'b0101001000: color_data = 12'b101100010010;
		10'b0101001001: color_data = 12'b101100010010;
		10'b0101001010: color_data = 12'b101100010010;
		10'b0101001011: color_data = 12'b101100010010;
		10'b0101001100: color_data = 12'b101100010010;
		10'b0101001101: color_data = 12'b101100010010;
		10'b0101001110: color_data = 12'b101100010010;
		10'b0101001111: color_data = 12'b101100010010;
		10'b0101010000: color_data = 12'b101100010010;
		10'b0101010001: color_data = 12'b101100010010;
		10'b0101010010: color_data = 12'b101100010010;
		10'b0101010011: color_data = 12'b101100010010;
		10'b0101010100: color_data = 12'b101100010010;
		10'b0101010101: color_data = 12'b101100100011;
		10'b0101010110: color_data = 12'b011011111110;
		10'b0101010111: color_data = 12'b011011111110;
		10'b0101100010: color_data = 12'b011011111110;
		10'b0101100011: color_data = 12'b011011111110;
		10'b0101100100: color_data = 12'b101100010010;
		10'b0101100101: color_data = 12'b101100010010;
		10'b0101100110: color_data = 12'b110000010010;
		10'b0101100111: color_data = 12'b101100010010;
		10'b0101101000: color_data = 12'b101100010010;
		10'b0101101001: color_data = 12'b101100010010;
		10'b0101101010: color_data = 12'b101100010010;
		10'b0101101011: color_data = 12'b101100010010;
		10'b0101101100: color_data = 12'b101100010010;
		10'b0101101101: color_data = 12'b101100010010;
		10'b0101101110: color_data = 12'b101100010010;
		10'b0101101111: color_data = 12'b101100010010;
		10'b0101110000: color_data = 12'b101100010010;
		10'b0101110001: color_data = 12'b101100010010;
		10'b0101110010: color_data = 12'b101100010010;
		10'b0101110011: color_data = 12'b101100010010;
		10'b0101110100: color_data = 12'b101100100011;
		10'b0101110101: color_data = 12'b101100010011;
		10'b0101110110: color_data = 12'b011011111110;
		10'b0101110111: color_data = 12'b011011111110;
		10'b0110000100: color_data = 12'b011011111110;
		10'b0110000101: color_data = 12'b011011111110;
		10'b0110000110: color_data = 12'b110000010011;
		10'b0110000111: color_data = 12'b101100010011;
		10'b0110001000: color_data = 12'b101100010010;
		10'b0110001001: color_data = 12'b101100010010;
		10'b0110001010: color_data = 12'b101100010010;
		10'b0110001011: color_data = 12'b101100010010;
		10'b0110001100: color_data = 12'b101100010010;
		10'b0110001101: color_data = 12'b101100010010;
		10'b0110001110: color_data = 12'b101100010010;
		10'b0110001111: color_data = 12'b101100010010;
		10'b0110010000: color_data = 12'b101100010010;
		10'b0110010001: color_data = 12'b110000010010;
		10'b0110010010: color_data = 12'b101100010010;
		10'b0110010011: color_data = 12'b110000010010;
		10'b0110010100: color_data = 12'b011011111110;
		10'b0110010101: color_data = 12'b011011111110;
		10'b0110100100: color_data = 12'b011011111110;
		10'b0110100101: color_data = 12'b011011111110;
		10'b0110100110: color_data = 12'b101100100010;
		10'b0110100111: color_data = 12'b101100100010;
		10'b0110101000: color_data = 12'b110000010010;
		10'b0110101001: color_data = 12'b101100010010;
		10'b0110101010: color_data = 12'b101100010010;
		10'b0110101011: color_data = 12'b101100010010;
		10'b0110101100: color_data = 12'b101100010010;
		10'b0110101101: color_data = 12'b101100010010;
		10'b0110101110: color_data = 12'b101100010010;
		10'b0110101111: color_data = 12'b101100010010;
		10'b0110110000: color_data = 12'b101100010010;
		10'b0110110001: color_data = 12'b101100010010;
		10'b0110110010: color_data = 12'b101100010010;
		10'b0110110011: color_data = 12'b101100100010;
		10'b0110110100: color_data = 12'b011011111110;
		10'b0110110101: color_data = 12'b011011111110;
		10'b0111000101: color_data = 12'b001000000000;
		10'b0111000110: color_data = 12'b011011111110;
		10'b0111000111: color_data = 12'b011011111110;
		10'b0111001000: color_data = 12'b101100010010;
		10'b0111001001: color_data = 12'b101100010010;
		10'b0111001010: color_data = 12'b101100010010;
		10'b0111001011: color_data = 12'b101100010010;
		10'b0111001100: color_data = 12'b101100010010;
		10'b0111001101: color_data = 12'b101100010010;
		10'b0111001110: color_data = 12'b101100010010;
		10'b0111001111: color_data = 12'b101100010010;
		10'b0111010000: color_data = 12'b101100010010;
		10'b0111010001: color_data = 12'b101100010011;
		10'b0111010010: color_data = 12'b011011111110;
		10'b0111010011: color_data = 12'b011011111110;
		10'b0111010100: color_data = 12'b000100000000;
		10'b0111100110: color_data = 12'b011011111110;
		10'b0111100111: color_data = 12'b011011111110;
		10'b0111101000: color_data = 12'b101100010010;
		10'b0111101001: color_data = 12'b101100010010;
		10'b0111101010: color_data = 12'b101100010010;
		10'b0111101011: color_data = 12'b101100010010;
		10'b0111101100: color_data = 12'b101100010010;
		10'b0111101101: color_data = 12'b101100010010;
		10'b0111101110: color_data = 12'b101100010010;
		10'b0111101111: color_data = 12'b101100010010;
		10'b0111110000: color_data = 12'b101100010010;
		10'b0111110001: color_data = 12'b110000010010;
		10'b0111110010: color_data = 12'b011011111110;
		10'b0111110011: color_data = 12'b011011111110;
		10'b1000001000: color_data = 12'b011011111110;
		10'b1000001001: color_data = 12'b011011111110;
		10'b1000001010: color_data = 12'b101100010010;
		10'b1000001011: color_data = 12'b101100010010;
		10'b1000001100: color_data = 12'b101100010010;
		10'b1000001101: color_data = 12'b101100010010;
		10'b1000001110: color_data = 12'b101100010011;
		10'b1000001111: color_data = 12'b110000010010;
		10'b1000010000: color_data = 12'b011011111110;
		10'b1000010001: color_data = 12'b011011111110;
		10'b1000101000: color_data = 12'b011011111110;
		10'b1000101001: color_data = 12'b011011111110;
		10'b1000101010: color_data = 12'b101100010010;
		10'b1000101011: color_data = 12'b101100010010;
		10'b1000101100: color_data = 12'b101100010010;
		10'b1000101101: color_data = 12'b101100010010;
		10'b1000101110: color_data = 12'b101100010011;
		10'b1000101111: color_data = 12'b101100010010;
		10'b1000110000: color_data = 12'b011011111110;
		10'b1000110001: color_data = 12'b011011111110;
		10'b1001001010: color_data = 12'b011011111110;
		10'b1001001011: color_data = 12'b011011111110;
		10'b1001001100: color_data = 12'b101100010010;
		10'b1001001101: color_data = 12'b101100100010;
		10'b1001001110: color_data = 12'b011011111110;
		10'b1001001111: color_data = 12'b011011111110;
		10'b1001101010: color_data = 12'b011011111110;
		10'b1001101011: color_data = 12'b011011111110;
		10'b1001101100: color_data = 12'b101100100010;
		10'b1001101101: color_data = 12'b101100010010;
		10'b1001101110: color_data = 12'b011011111110;
		10'b1001101111: color_data = 12'b011011111110;
		10'b1010001010: color_data = 12'b011011111110;
		10'b1010001011: color_data = 12'b011011111110;
		10'b1010001100: color_data = 12'b110000010010;
		10'b1010001101: color_data = 12'b101100010010;
		10'b1010001110: color_data = 12'b011011111110;
		10'b1010001111: color_data = 12'b011011111110;
		10'b1010101100: color_data = 12'b011011111110;
		10'b1010101101: color_data = 12'b011011111110;
		10'b1011001100: color_data = 12'b011011111110;
		10'b1011001101: color_data = 12'b011011111110;
		default: color_data = 12'b000000000000;
	endcase
endmodule