`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.01.2025 15:05:54
// Design Name: 
// Module Name: player_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

	module player_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: color_data = 12'b111100010001;
		12'b000000000001: color_data = 12'b111100010001;
		12'b000000000010: color_data = 12'b111100010001;
		12'b000000000011: color_data = 12'b111100010001;
		12'b000000000100: color_data = 12'b111100010001;
		12'b000000000101: color_data = 12'b111100010001;
		12'b000000000110: color_data = 12'b111100010001;
		12'b000000000111: color_data = 12'b111100010001;
		12'b000000001000: color_data = 12'b111100010001;
		12'b000000001001: color_data = 12'b111100010001;
		12'b000000001010: color_data = 12'b111100010001;
		12'b000000001011: color_data = 12'b111100010001;
		12'b000000001100: color_data = 12'b111100010001;
		12'b000000001101: color_data = 12'b111100010001;
		12'b000000010001: color_data = 12'b111100010001;
		12'b000000010010: color_data = 12'b111100010001;
		12'b000000010011: color_data = 12'b111100010001;
		12'b000000010100: color_data = 12'b111100010001;
		12'b000010000000: color_data = 12'b111100010001;
		12'b000010000001: color_data = 12'b111100010001;
		12'b000010000010: color_data = 12'b111100010001;
		12'b000010000011: color_data = 12'b111100010001;
		12'b000010000100: color_data = 12'b111100010001;
		12'b000010000101: color_data = 12'b111100010001;
		12'b000010000110: color_data = 12'b111100010001;
		12'b000010000111: color_data = 12'b111100010001;
		12'b000010001000: color_data = 12'b111100010001;
		12'b000010001001: color_data = 12'b111100010001;
		12'b000010001010: color_data = 12'b111100010001;
		12'b000010001011: color_data = 12'b111100010001;
		12'b000010001100: color_data = 12'b111100010001;
		12'b000010001101: color_data = 12'b111100010001;
		12'b000010010001: color_data = 12'b111100010001;
		12'b000010010010: color_data = 12'b111100010001;
		12'b000010010011: color_data = 12'b111100010001;
		12'b000010010100: color_data = 12'b111100010001;
		12'b000100000000: color_data = 12'b111100010001;
		12'b000100000001: color_data = 12'b111100010001;
		12'b000100000010: color_data = 12'b111100010001;
		12'b000100000011: color_data = 12'b111100010001;
		12'b000100000100: color_data = 12'b111100010001;
		12'b000100000101: color_data = 12'b111100010001;
		12'b000100000110: color_data = 12'b111100010001;
		12'b000100000111: color_data = 12'b111100010001;
		12'b000100001000: color_data = 12'b111100010001;
		12'b000100001001: color_data = 12'b111100010001;
		12'b000100001010: color_data = 12'b111100010001;
		12'b000100001011: color_data = 12'b111100010001;
		12'b000100001100: color_data = 12'b111100010001;
		12'b000100001101: color_data = 12'b111100010001;
		12'b000100010001: color_data = 12'b111100010001;
		12'b000100010010: color_data = 12'b111100010001;
		12'b000100010011: color_data = 12'b111100010001;
		12'b000100010100: color_data = 12'b111100010001;
		12'b000110000000: color_data = 12'b111100010001;
		12'b000110000001: color_data = 12'b111100010001;
		12'b000110000010: color_data = 12'b111100010001;
		12'b000110000011: color_data = 12'b111100010001;
		12'b000110001011: color_data = 12'b111100010001;
		12'b000110001100: color_data = 12'b111100010001;
		12'b000110001101: color_data = 12'b111100010001;
		12'b000110010001: color_data = 12'b111100010001;
		12'b000110010010: color_data = 12'b111100010001;
		12'b000110010011: color_data = 12'b111100010001;
		12'b000110010100: color_data = 12'b111100010001;
		12'b001000000000: color_data = 12'b111100010001;
		12'b001000000001: color_data = 12'b111100010001;
		12'b001000000010: color_data = 12'b111100010001;
		12'b001000000011: color_data = 12'b111100010001;
		12'b001000001011: color_data = 12'b111100010001;
		12'b001000001100: color_data = 12'b111100010001;
		12'b001000001101: color_data = 12'b111100010001;
		12'b001000010001: color_data = 12'b111100010001;
		12'b001000010010: color_data = 12'b111100010001;
		12'b001000010011: color_data = 12'b111100010001;
		12'b001000010100: color_data = 12'b111100010001;
		12'b001010000000: color_data = 12'b111100010001;
		12'b001010000001: color_data = 12'b111100010001;
		12'b001010000010: color_data = 12'b111100010001;
		12'b001010000011: color_data = 12'b111100010001;
		12'b001010001011: color_data = 12'b111100010001;
		12'b001010001100: color_data = 12'b111100010001;
		12'b001010001101: color_data = 12'b111100010001;
		12'b001010010001: color_data = 12'b111100010001;
		12'b001010010010: color_data = 12'b111100010001;
		12'b001010010011: color_data = 12'b111100010001;
		12'b001010010100: color_data = 12'b111100010001;
		12'b001100000000: color_data = 12'b111100010001;
		12'b001100000001: color_data = 12'b111100010001;
		12'b001100000010: color_data = 12'b111100010001;
		12'b001100000011: color_data = 12'b111100010001;
		12'b001100000100: color_data = 12'b111100010001;
		12'b001100000101: color_data = 12'b111100010001;
		12'b001100000110: color_data = 12'b111100010001;
		12'b001100000111: color_data = 12'b111100010001;
		12'b001100001000: color_data = 12'b111100010001;
		12'b001100001001: color_data = 12'b111100010001;
		12'b001100001010: color_data = 12'b111100010001;
		12'b001100001011: color_data = 12'b111100010001;
		12'b001100001100: color_data = 12'b111100010001;
		12'b001100001101: color_data = 12'b111100010001;
		12'b001100010001: color_data = 12'b111100010001;
		12'b001100010010: color_data = 12'b111100010001;
		12'b001100010011: color_data = 12'b111100010001;
		12'b001100010100: color_data = 12'b111100010001;
		12'b001100011100: color_data = 12'b111100010001;
		12'b001100011101: color_data = 12'b111100010001;
		12'b001100011110: color_data = 12'b111100010001;
		12'b001100011111: color_data = 12'b111100010001;
		12'b001100100000: color_data = 12'b111100010001;
		12'b001100100001: color_data = 12'b111100010001;
		12'b001100100110: color_data = 12'b111100010001;
		12'b001100100111: color_data = 12'b111100010001;
		12'b001100101000: color_data = 12'b111100010001;
		12'b001100101100: color_data = 12'b111100010001;
		12'b001100101101: color_data = 12'b111100010001;
		12'b001100101110: color_data = 12'b111100010001;
		12'b001100101111: color_data = 12'b111100010001;
		12'b001100110011: color_data = 12'b111100010001;
		12'b001100110100: color_data = 12'b111100010001;
		12'b001100110101: color_data = 12'b111100010001;
		12'b001100110110: color_data = 12'b111100010001;
		12'b001100110111: color_data = 12'b111100010001;
		12'b001100111000: color_data = 12'b111100010001;
		12'b001100111001: color_data = 12'b111100010001;
		12'b001100111010: color_data = 12'b111100010001;
		12'b001100111011: color_data = 12'b111100010001;
		12'b001100111100: color_data = 12'b111100010001;
		12'b001101000001: color_data = 12'b111100010001;
		12'b001101000010: color_data = 12'b111100010001;
		12'b001101000011: color_data = 12'b111100010001;
		12'b001101000100: color_data = 12'b111100010001;
		12'b001101000101: color_data = 12'b111100010001;
		12'b001101000110: color_data = 12'b111100010001;
		12'b001110000000: color_data = 12'b111100010001;
		12'b001110000001: color_data = 12'b111100010001;
		12'b001110000010: color_data = 12'b111100010001;
		12'b001110000011: color_data = 12'b111100010001;
		12'b001110000100: color_data = 12'b111100010001;
		12'b001110000101: color_data = 12'b111100010001;
		12'b001110000110: color_data = 12'b111100010001;
		12'b001110000111: color_data = 12'b111100010001;
		12'b001110001000: color_data = 12'b111100010001;
		12'b001110001001: color_data = 12'b111100010001;
		12'b001110001010: color_data = 12'b111100010001;
		12'b001110001011: color_data = 12'b111100010001;
		12'b001110001100: color_data = 12'b111100010001;
		12'b001110001101: color_data = 12'b111100010001;
		12'b001110010001: color_data = 12'b111100010001;
		12'b001110010010: color_data = 12'b111100010001;
		12'b001110010011: color_data = 12'b111100010001;
		12'b001110010100: color_data = 12'b111100010001;
		12'b001110011100: color_data = 12'b111100010001;
		12'b001110011101: color_data = 12'b111100010001;
		12'b001110011110: color_data = 12'b111100010001;
		12'b001110011111: color_data = 12'b111100010001;
		12'b001110100000: color_data = 12'b111100010001;
		12'b001110100001: color_data = 12'b111100010001;
		12'b001110100110: color_data = 12'b111100010001;
		12'b001110100111: color_data = 12'b111100010001;
		12'b001110101000: color_data = 12'b111100010001;
		12'b001110101100: color_data = 12'b111100010001;
		12'b001110101101: color_data = 12'b111100010001;
		12'b001110101110: color_data = 12'b111100010001;
		12'b001110101111: color_data = 12'b111100010001;
		12'b001110110011: color_data = 12'b111100010001;
		12'b001110110100: color_data = 12'b111100010001;
		12'b001110110101: color_data = 12'b111100010001;
		12'b001110110110: color_data = 12'b111100010001;
		12'b001110110111: color_data = 12'b111100010001;
		12'b001110111000: color_data = 12'b111100010001;
		12'b001110111001: color_data = 12'b111100010001;
		12'b001110111010: color_data = 12'b111100010001;
		12'b001110111011: color_data = 12'b111100010001;
		12'b001110111100: color_data = 12'b111100010001;
		12'b001111000001: color_data = 12'b111100010001;
		12'b001111000010: color_data = 12'b111100010001;
		12'b001111000011: color_data = 12'b111100010001;
		12'b001111000100: color_data = 12'b111100010001;
		12'b001111000101: color_data = 12'b111100010001;
		12'b001111000110: color_data = 12'b111100010001;
		12'b010000000000: color_data = 12'b111100010001;
		12'b010000000001: color_data = 12'b111100010001;
		12'b010000000010: color_data = 12'b111100010001;
		12'b010000000011: color_data = 12'b111100010001;
		12'b010000000100: color_data = 12'b111100010001;
		12'b010000000101: color_data = 12'b111100010001;
		12'b010000000110: color_data = 12'b111100010001;
		12'b010000000111: color_data = 12'b111100010001;
		12'b010000001000: color_data = 12'b111100010001;
		12'b010000001001: color_data = 12'b111100010001;
		12'b010000001010: color_data = 12'b111100010001;
		12'b010000001011: color_data = 12'b111100010001;
		12'b010000001100: color_data = 12'b111100010001;
		12'b010000001101: color_data = 12'b111100010001;
		12'b010000010001: color_data = 12'b111100010001;
		12'b010000010010: color_data = 12'b111100010001;
		12'b010000010011: color_data = 12'b111100010001;
		12'b010000010100: color_data = 12'b111100010001;
		12'b010000011100: color_data = 12'b111100010001;
		12'b010000011101: color_data = 12'b111100010001;
		12'b010000011110: color_data = 12'b111100010001;
		12'b010000011111: color_data = 12'b111100010001;
		12'b010000100000: color_data = 12'b111100010001;
		12'b010000100001: color_data = 12'b111100010001;
		12'b010000100110: color_data = 12'b111100010001;
		12'b010000100111: color_data = 12'b111100010001;
		12'b010000101000: color_data = 12'b111100010001;
		12'b010000101100: color_data = 12'b111100010001;
		12'b010000101101: color_data = 12'b111100010001;
		12'b010000101110: color_data = 12'b111100010001;
		12'b010000101111: color_data = 12'b111100010001;
		12'b010000110011: color_data = 12'b111100010001;
		12'b010000110100: color_data = 12'b111100010001;
		12'b010000110101: color_data = 12'b111100010001;
		12'b010000110110: color_data = 12'b111100010001;
		12'b010000110111: color_data = 12'b111100010001;
		12'b010000111000: color_data = 12'b111100010001;
		12'b010000111001: color_data = 12'b111100010001;
		12'b010000111010: color_data = 12'b111100010001;
		12'b010000111011: color_data = 12'b111100010001;
		12'b010000111100: color_data = 12'b111100010001;
		12'b010001000001: color_data = 12'b111100010001;
		12'b010001000010: color_data = 12'b111100010001;
		12'b010001000011: color_data = 12'b111100010001;
		12'b010001000100: color_data = 12'b111100010001;
		12'b010001000101: color_data = 12'b111100010001;
		12'b010001000110: color_data = 12'b111100010001;
		12'b010010000000: color_data = 12'b111100010001;
		12'b010010000001: color_data = 12'b111100010001;
		12'b010010000010: color_data = 12'b111100010001;
		12'b010010000011: color_data = 12'b111100010001;
		12'b010010010001: color_data = 12'b111100010001;
		12'b010010010010: color_data = 12'b111100010001;
		12'b010010010011: color_data = 12'b111100010001;
		12'b010010010100: color_data = 12'b111100010001;
		12'b010010011000: color_data = 12'b111100010001;
		12'b010010011001: color_data = 12'b111100010001;
		12'b010010011010: color_data = 12'b111100010001;
		12'b010010011011: color_data = 12'b111100010001;
		12'b010010011111: color_data = 12'b111100010001;
		12'b010010100000: color_data = 12'b111100010001;
		12'b010010100001: color_data = 12'b111100010001;
		12'b010010100110: color_data = 12'b111100010001;
		12'b010010100111: color_data = 12'b111100010001;
		12'b010010101000: color_data = 12'b111100010001;
		12'b010010101100: color_data = 12'b111100010001;
		12'b010010101101: color_data = 12'b111100010001;
		12'b010010101110: color_data = 12'b111100010001;
		12'b010010101111: color_data = 12'b111100010001;
		12'b010010110011: color_data = 12'b111100010001;
		12'b010010110100: color_data = 12'b111100010001;
		12'b010010110101: color_data = 12'b111100010001;
		12'b010010110110: color_data = 12'b111100010001;
		12'b010010111010: color_data = 12'b111100010001;
		12'b010010111011: color_data = 12'b111100010001;
		12'b010010111100: color_data = 12'b111100010001;
		12'b010011000001: color_data = 12'b111100010001;
		12'b010011000010: color_data = 12'b111100010001;
		12'b010011000011: color_data = 12'b111100010001;
		12'b010100000000: color_data = 12'b111100010001;
		12'b010100000001: color_data = 12'b111100010001;
		12'b010100000010: color_data = 12'b111100010001;
		12'b010100000011: color_data = 12'b111100010001;
		12'b010100010001: color_data = 12'b111100010001;
		12'b010100010010: color_data = 12'b111100010001;
		12'b010100010011: color_data = 12'b111100010001;
		12'b010100010100: color_data = 12'b111100010001;
		12'b010100011000: color_data = 12'b111100010001;
		12'b010100011001: color_data = 12'b111100010001;
		12'b010100011010: color_data = 12'b111100010001;
		12'b010100011011: color_data = 12'b111100010001;
		12'b010100011111: color_data = 12'b111100010001;
		12'b010100100000: color_data = 12'b111100010001;
		12'b010100100001: color_data = 12'b111100010001;
		12'b010100100110: color_data = 12'b111100010001;
		12'b010100100111: color_data = 12'b111100010001;
		12'b010100101000: color_data = 12'b111100010001;
		12'b010100101100: color_data = 12'b111100010001;
		12'b010100101101: color_data = 12'b111100010001;
		12'b010100101110: color_data = 12'b111100010001;
		12'b010100101111: color_data = 12'b111100010001;
		12'b010100110011: color_data = 12'b111100010001;
		12'b010100110100: color_data = 12'b111100010001;
		12'b010100110101: color_data = 12'b111100010001;
		12'b010100110110: color_data = 12'b111100010001;
		12'b010100111010: color_data = 12'b111100010001;
		12'b010100111011: color_data = 12'b111100010001;
		12'b010100111100: color_data = 12'b111100010001;
		12'b010101000001: color_data = 12'b111100010001;
		12'b010101000010: color_data = 12'b111100010001;
		12'b010101000011: color_data = 12'b111100010001;
		12'b010110000000: color_data = 12'b111100010001;
		12'b010110000001: color_data = 12'b111100010001;
		12'b010110000010: color_data = 12'b111100010001;
		12'b010110000011: color_data = 12'b111100010001;
		12'b010110010001: color_data = 12'b111100010001;
		12'b010110010010: color_data = 12'b111100010001;
		12'b010110010011: color_data = 12'b111100010001;
		12'b010110010100: color_data = 12'b111100010001;
		12'b010110011000: color_data = 12'b111100010001;
		12'b010110011001: color_data = 12'b111100010001;
		12'b010110011010: color_data = 12'b111100010001;
		12'b010110011011: color_data = 12'b111100010001;
		12'b010110011111: color_data = 12'b111100010001;
		12'b010110100000: color_data = 12'b111100010001;
		12'b010110100001: color_data = 12'b111100010001;
		12'b010110100110: color_data = 12'b111100010001;
		12'b010110100111: color_data = 12'b111100010001;
		12'b010110101000: color_data = 12'b111100010001;
		12'b010110101100: color_data = 12'b111100010001;
		12'b010110101101: color_data = 12'b111100010001;
		12'b010110101110: color_data = 12'b111100010001;
		12'b010110101111: color_data = 12'b111100010001;
		12'b010110110011: color_data = 12'b111100010001;
		12'b010110110100: color_data = 12'b111100010001;
		12'b010110110101: color_data = 12'b111100010001;
		12'b010110110110: color_data = 12'b111100010001;
		12'b010110111010: color_data = 12'b111100010001;
		12'b010110111011: color_data = 12'b111100010001;
		12'b010110111100: color_data = 12'b111100010001;
		12'b010111000001: color_data = 12'b111100010001;
		12'b010111000010: color_data = 12'b111100010001;
		12'b010111000011: color_data = 12'b111100010001;
		12'b011000000000: color_data = 12'b111100010001;
		12'b011000000001: color_data = 12'b111100010001;
		12'b011000000010: color_data = 12'b111100010001;
		12'b011000000011: color_data = 12'b111100010001;
		12'b011000010001: color_data = 12'b111100010001;
		12'b011000010010: color_data = 12'b111100010001;
		12'b011000010011: color_data = 12'b111100010001;
		12'b011000010100: color_data = 12'b111100010001;
		12'b011000011000: color_data = 12'b111100010001;
		12'b011000011001: color_data = 12'b111100010001;
		12'b011000011010: color_data = 12'b111100010001;
		12'b011000011011: color_data = 12'b111100010001;
		12'b011000011100: color_data = 12'b111100010001;
		12'b011000011101: color_data = 12'b111100010001;
		12'b011000011110: color_data = 12'b111100010001;
		12'b011000011111: color_data = 12'b111100010001;
		12'b011000100000: color_data = 12'b111100010001;
		12'b011000100001: color_data = 12'b111100010001;
		12'b011000100110: color_data = 12'b111100010001;
		12'b011000100111: color_data = 12'b111100010001;
		12'b011000101000: color_data = 12'b111100010001;
		12'b011000101001: color_data = 12'b111100010001;
		12'b011000101010: color_data = 12'b111100010001;
		12'b011000101011: color_data = 12'b111100010001;
		12'b011000101100: color_data = 12'b111100010001;
		12'b011000101101: color_data = 12'b111100010001;
		12'b011000101110: color_data = 12'b111100010001;
		12'b011000101111: color_data = 12'b111100010001;
		12'b011000110011: color_data = 12'b111100010001;
		12'b011000110100: color_data = 12'b111100010001;
		12'b011000110101: color_data = 12'b111100010001;
		12'b011000110110: color_data = 12'b111100010001;
		12'b011000110111: color_data = 12'b111100010001;
		12'b011000111000: color_data = 12'b111100010001;
		12'b011000111001: color_data = 12'b111100010001;
		12'b011001000001: color_data = 12'b111100010001;
		12'b011001000010: color_data = 12'b111100010001;
		12'b011001000011: color_data = 12'b111100010001;
		12'b011010000000: color_data = 12'b111100010001;
		12'b011010000001: color_data = 12'b111100010001;
		12'b011010000010: color_data = 12'b111100010001;
		12'b011010000011: color_data = 12'b111100010001;
		12'b011010010001: color_data = 12'b111100010001;
		12'b011010010010: color_data = 12'b111100010001;
		12'b011010010011: color_data = 12'b111100010001;
		12'b011010010100: color_data = 12'b111100010001;
		12'b011010011000: color_data = 12'b111100010001;
		12'b011010011001: color_data = 12'b111100010001;
		12'b011010011010: color_data = 12'b111100010001;
		12'b011010011011: color_data = 12'b111100010001;
		12'b011010011100: color_data = 12'b111100010001;
		12'b011010011101: color_data = 12'b111100010001;
		12'b011010011110: color_data = 12'b111100010001;
		12'b011010011111: color_data = 12'b111100010001;
		12'b011010100000: color_data = 12'b111100010001;
		12'b011010100001: color_data = 12'b111100010001;
		12'b011010100110: color_data = 12'b111100010001;
		12'b011010100111: color_data = 12'b111100010001;
		12'b011010101000: color_data = 12'b111100010001;
		12'b011010101001: color_data = 12'b111100010001;
		12'b011010101010: color_data = 12'b111100010001;
		12'b011010101011: color_data = 12'b111100010001;
		12'b011010101100: color_data = 12'b111100010001;
		12'b011010101101: color_data = 12'b111100010001;
		12'b011010101110: color_data = 12'b111100010001;
		12'b011010101111: color_data = 12'b111100010001;
		12'b011010110011: color_data = 12'b111100010001;
		12'b011010110100: color_data = 12'b111100010001;
		12'b011010110101: color_data = 12'b111100010001;
		12'b011010110110: color_data = 12'b111100010001;
		12'b011010110111: color_data = 12'b111100010001;
		12'b011010111000: color_data = 12'b111100010001;
		12'b011010111001: color_data = 12'b111100010001;
		12'b011011000001: color_data = 12'b111100010001;
		12'b011011000010: color_data = 12'b111100010001;
		12'b011011000011: color_data = 12'b111100010001;
		12'b011100000000: color_data = 12'b111100010001;
		12'b011100000001: color_data = 12'b111100010001;
		12'b011100000010: color_data = 12'b111100010001;
		12'b011100000011: color_data = 12'b111100010001;
		12'b011100010001: color_data = 12'b111100010001;
		12'b011100010010: color_data = 12'b111100010001;
		12'b011100010011: color_data = 12'b111100010001;
		12'b011100010100: color_data = 12'b111100010001;
		12'b011100011000: color_data = 12'b111100010001;
		12'b011100011001: color_data = 12'b111100010001;
		12'b011100011010: color_data = 12'b111100010001;
		12'b011100011011: color_data = 12'b111100010001;
		12'b011100011100: color_data = 12'b111100010001;
		12'b011100011101: color_data = 12'b111100010001;
		12'b011100011110: color_data = 12'b111100010001;
		12'b011100011111: color_data = 12'b111100010001;
		12'b011100100000: color_data = 12'b111100010001;
		12'b011100100001: color_data = 12'b111100010001;
		12'b011100100110: color_data = 12'b111100010001;
		12'b011100100111: color_data = 12'b111100010001;
		12'b011100101000: color_data = 12'b111100010001;
		12'b011100101001: color_data = 12'b111100010001;
		12'b011100101010: color_data = 12'b111100010001;
		12'b011100101011: color_data = 12'b111100010001;
		12'b011100101100: color_data = 12'b111100010001;
		12'b011100101101: color_data = 12'b111100010001;
		12'b011100101110: color_data = 12'b111100010001;
		12'b011100101111: color_data = 12'b111100010001;
		12'b011100110011: color_data = 12'b111100010001;
		12'b011100110100: color_data = 12'b111100010001;
		12'b011100110101: color_data = 12'b111100010001;
		12'b011100110110: color_data = 12'b111100010001;
		12'b011100110111: color_data = 12'b111100010001;
		12'b011100111000: color_data = 12'b111100010001;
		12'b011100111001: color_data = 12'b111100010001;
		12'b011101000001: color_data = 12'b111100010001;
		12'b011101000010: color_data = 12'b111100010001;
		12'b011101000011: color_data = 12'b111100010001;
		12'b011110101100: color_data = 12'b111100010001;
		12'b011110101101: color_data = 12'b111100010001;
		12'b011110101110: color_data = 12'b111100010001;
		12'b011110101111: color_data = 12'b111100010001;
		12'b100000101100: color_data = 12'b111100010001;
		12'b100000101101: color_data = 12'b111100010001;
		12'b100000101110: color_data = 12'b111100010001;
		12'b100000101111: color_data = 12'b111100010001;
		12'b100010101100: color_data = 12'b111100010001;
		12'b100010101101: color_data = 12'b111100010001;
		12'b100010101110: color_data = 12'b111100010001;
		12'b100010101111: color_data = 12'b111100010001;
		12'b100100100110: color_data = 12'b111100010001;
		12'b100100100111: color_data = 12'b111100010001;
		12'b100100101000: color_data = 12'b111100010001;
		12'b100100101001: color_data = 12'b111100010001;
		12'b100100101010: color_data = 12'b111100010001;
		12'b100100101011: color_data = 12'b111100010001;
		12'b100100101100: color_data = 12'b111100010001;
		12'b100100101101: color_data = 12'b111100010001;
		12'b100100101110: color_data = 12'b111100010001;
		12'b100100101111: color_data = 12'b111100010001;
		12'b100110100110: color_data = 12'b111100010001;
		12'b100110100111: color_data = 12'b111100010001;
		12'b100110101000: color_data = 12'b111100010001;
		12'b100110101001: color_data = 12'b111100010001;
		12'b100110101010: color_data = 12'b111100010001;
		12'b100110101011: color_data = 12'b111100010001;
		12'b100110101100: color_data = 12'b111100010001;
		12'b100110101101: color_data = 12'b111100010001;
		12'b100110101110: color_data = 12'b111100010001;
		12'b100110101111: color_data = 12'b111100010001;
		12'b101000100110: color_data = 12'b111100010001;
		12'b101000100111: color_data = 12'b111100010001;
		12'b101000101000: color_data = 12'b111100010001;
		12'b101000101001: color_data = 12'b111100010001;
		12'b101000101010: color_data = 12'b111100010001;
		12'b101000101011: color_data = 12'b111100010001;
		12'b101000101100: color_data = 12'b111100010001;
		12'b101000101101: color_data = 12'b111100010001;
		12'b101000101110: color_data = 12'b111100010001;
		12'b101000101111: color_data = 12'b111100010001;
		default: color_data = 12'b000000000000;
	endcase
endmodule
