module top(

);
