		module yes_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		11'b00000000000: color_data = 12'b110011110111;
		11'b00000000001: color_data = 12'b110011110111;
		11'b00000000010: color_data = 12'b110011110111;
		11'b00000001000: color_data = 12'b110011110111;
		11'b00000001001: color_data = 12'b110011110111;
		11'b00000001010: color_data = 12'b110011110111;
		11'b00001000000: color_data = 12'b110011110111;
		11'b00001000001: color_data = 12'b110011110111;
		11'b00001000010: color_data = 12'b110011110111;
		11'b00001000011: color_data = 12'b110011110111;
		11'b00001000111: color_data = 12'b110011110111;
		11'b00001001000: color_data = 12'b110011110111;
		11'b00001001001: color_data = 12'b110011110111;
		11'b00001001101: color_data = 12'b110011110111;
		11'b00001001110: color_data = 12'b110011110111;
		11'b00001001111: color_data = 12'b110011110111;
		11'b00001010000: color_data = 12'b110011110111;
		11'b00001010001: color_data = 12'b110011110111;
		11'b00001010010: color_data = 12'b110011110111;
		11'b00001010011: color_data = 12'b110011110111;
		11'b00001010100: color_data = 12'b110011110111;
		11'b00001010101: color_data = 12'b110011110111;
		11'b00001010110: color_data = 12'b110011110111;
		11'b00001011010: color_data = 12'b110011110111;
		11'b00001011011: color_data = 12'b110011110111;
		11'b00001011100: color_data = 12'b110011110111;
		11'b00001011101: color_data = 12'b110011110111;
		11'b00001011110: color_data = 12'b110011110111;
		11'b00001011111: color_data = 12'b110011110111;
		11'b00001100000: color_data = 12'b110011110111;
		11'b00001100001: color_data = 12'b110011110111;
		11'b00001100010: color_data = 12'b110011110111;
		11'b00010000000: color_data = 12'b110011110111;
		11'b00010000001: color_data = 12'b110011110111;
		11'b00010000010: color_data = 12'b110011110111;
		11'b00010000011: color_data = 12'b110011110111;
		11'b00010000111: color_data = 12'b110011110111;
		11'b00010001000: color_data = 12'b110011110111;
		11'b00010001001: color_data = 12'b110011110111;
		11'b00010001101: color_data = 12'b110011110111;
		11'b00010001110: color_data = 12'b110011110111;
		11'b00010001111: color_data = 12'b110011110111;
		11'b00010010101: color_data = 12'b110011110111;
		11'b00010010110: color_data = 12'b110011110111;
		11'b00010010111: color_data = 12'b110011110111;
		11'b00010011010: color_data = 12'b110011110111;
		11'b00010011011: color_data = 12'b110011110111;
		11'b00010100010: color_data = 12'b110011110111;
		11'b00010100011: color_data = 12'b110011110111;
		11'b00011000001: color_data = 12'b110011110111;
		11'b00011000010: color_data = 12'b110011110111;
		11'b00011000100: color_data = 12'b110011110111;
		11'b00011000111: color_data = 12'b110011110111;
		11'b00011001000: color_data = 12'b110011110111;
		11'b00011001010: color_data = 12'b110011110111;
		11'b00011001101: color_data = 12'b110011110111;
		11'b00011001110: color_data = 12'b110011110111;
		11'b00011001111: color_data = 12'b110011110111;
		11'b00011010110: color_data = 12'b110011110111;
		11'b00011010111: color_data = 12'b110011110111;
		11'b00011011001: color_data = 12'b110011110111;
		11'b00011011010: color_data = 12'b110011110111;
		11'b00011011011: color_data = 12'b110011110111;
		11'b00011100010: color_data = 12'b110011110111;
		11'b00011100011: color_data = 12'b110011110111;
		11'b00011100100: color_data = 12'b110011110111;
		11'b00100000010: color_data = 12'b110011110111;
		11'b00100000011: color_data = 12'b110011110111;
		11'b00100000101: color_data = 12'b110011110111;
		11'b00100000111: color_data = 12'b110011110111;
		11'b00100001000: color_data = 12'b110011110111;
		11'b00100001010: color_data = 12'b110011110111;
		11'b00100001101: color_data = 12'b110011110111;
		11'b00100001110: color_data = 12'b110011110111;
		11'b00100001111: color_data = 12'b110011110111;
		11'b00100011001: color_data = 12'b110011110111;
		11'b00100011011: color_data = 12'b110011110111;
		11'b00100100100: color_data = 12'b110011110111;
		11'b00101000010: color_data = 12'b110011110111;
		11'b00101000011: color_data = 12'b110011110111;
		11'b00101000101: color_data = 12'b110011110111;
		11'b00101000110: color_data = 12'b110011110111;
		11'b00101000111: color_data = 12'b110011110111;
		11'b00101001001: color_data = 12'b110011110111;
		11'b00101001101: color_data = 12'b110011110111;
		11'b00101001110: color_data = 12'b110011110111;
		11'b00101001111: color_data = 12'b110011110111;
		11'b00101011001: color_data = 12'b110011110111;
		11'b00101011011: color_data = 12'b110011110111;
		11'b00110000011: color_data = 12'b110011110111;
		11'b00110000100: color_data = 12'b110011110111;
		11'b00110000101: color_data = 12'b110011110111;
		11'b00110000110: color_data = 12'b110011110111;
		11'b00110000111: color_data = 12'b110011110111;
		11'b00110001001: color_data = 12'b110011110111;
		11'b00110001101: color_data = 12'b110011110111;
		11'b00110001110: color_data = 12'b110011110111;
		11'b00110001111: color_data = 12'b110011110111;
		11'b00110011001: color_data = 12'b110011110111;
		11'b00110011011: color_data = 12'b110011110111;
		11'b00111000011: color_data = 12'b110011110111;
		11'b00111000100: color_data = 12'b110011110111;
		11'b00111000101: color_data = 12'b110011110111;
		11'b00111000110: color_data = 12'b110011110111;
		11'b00111001000: color_data = 12'b110011110111;
		11'b00111001101: color_data = 12'b110011110111;
		11'b00111001110: color_data = 12'b110011110111;
		11'b00111001111: color_data = 12'b110011110111;
		11'b00111011001: color_data = 12'b110011110111;
		11'b00111011010: color_data = 12'b110011110111;
		11'b00111011011: color_data = 12'b110011110111;
		11'b01000000011: color_data = 12'b110011110111;
		11'b01000000100: color_data = 12'b110011110111;
		11'b01000000101: color_data = 12'b110011110111;
		11'b01000000110: color_data = 12'b110011110111;
		11'b01000001000: color_data = 12'b110011110111;
		11'b01000001101: color_data = 12'b110011110111;
		11'b01000001110: color_data = 12'b110011110111;
		11'b01000001111: color_data = 12'b110011110111;
		11'b01000010000: color_data = 12'b110011110111;
		11'b01000010001: color_data = 12'b110011110111;
		11'b01000010010: color_data = 12'b110011110111;
		11'b01000010011: color_data = 12'b110011110111;
		11'b01000010100: color_data = 12'b110011110111;
		11'b01000010101: color_data = 12'b110011110111;
		11'b01000011010: color_data = 12'b110011110111;
		11'b01000011011: color_data = 12'b110011110111;
		11'b01000011100: color_data = 12'b110011110111;
		11'b01000011101: color_data = 12'b110011110111;
		11'b01000011110: color_data = 12'b110011110111;
		11'b01000011111: color_data = 12'b110011110111;
		11'b01000100000: color_data = 12'b110011110111;
		11'b01000100001: color_data = 12'b110011110111;
		11'b01001000100: color_data = 12'b110011110111;
		11'b01001000101: color_data = 12'b110011110111;
		11'b01001000110: color_data = 12'b110011110111;
		11'b01001000111: color_data = 12'b110011110111;
		11'b01001001101: color_data = 12'b110011110111;
		11'b01001001110: color_data = 12'b110011110111;
		11'b01001001111: color_data = 12'b110011110111;
		11'b01001010000: color_data = 12'b110011110111;
		11'b01001010001: color_data = 12'b110011110111;
		11'b01001010010: color_data = 12'b110011110111;
		11'b01001010011: color_data = 12'b110011110111;
		11'b01001010100: color_data = 12'b110011110111;
		11'b01001010101: color_data = 12'b110011110111;
		11'b01001011010: color_data = 12'b110011110111;
		11'b01001011011: color_data = 12'b110011110111;
		11'b01001011100: color_data = 12'b110011110111;
		11'b01001011101: color_data = 12'b110011110111;
		11'b01001011110: color_data = 12'b110011110111;
		11'b01001011111: color_data = 12'b110011110111;
		11'b01001100000: color_data = 12'b110011110111;
		11'b01001100001: color_data = 12'b110011110111;
		11'b01001100010: color_data = 12'b110011110111;
		11'b01010000100: color_data = 12'b110011110111;
		11'b01010000101: color_data = 12'b110011110111;
		11'b01010000110: color_data = 12'b110011110111;
		11'b01010000111: color_data = 12'b110011110111;
		11'b01010001101: color_data = 12'b110011110111;
		11'b01010001110: color_data = 12'b110011110111;
		11'b01010001111: color_data = 12'b110011110111;
		11'b01010100010: color_data = 12'b110011110111;
		11'b01010100011: color_data = 12'b110011110111;
		11'b01010100100: color_data = 12'b110011110111;
		11'b01011000100: color_data = 12'b110011110111;
		11'b01011000101: color_data = 12'b110011110111;
		11'b01011000110: color_data = 12'b110011110111;
		11'b01011000111: color_data = 12'b110011110111;
		11'b01011001101: color_data = 12'b110011110111;
		11'b01011001110: color_data = 12'b110011110111;
		11'b01011001111: color_data = 12'b110011110111;
		11'b01011100011: color_data = 12'b110011110111;
		11'b01011100100: color_data = 12'b110011110111;
		11'b01100000100: color_data = 12'b110011110111;
		11'b01100000101: color_data = 12'b110011110111;
		11'b01100000110: color_data = 12'b110011110111;
		11'b01100000111: color_data = 12'b110011110111;
		11'b01100001101: color_data = 12'b110011110111;
		11'b01100001110: color_data = 12'b110011110111;
		11'b01100001111: color_data = 12'b110011110111;
		11'b01100100011: color_data = 12'b110011110111;
		11'b01100100100: color_data = 12'b110011110111;
		11'b01101000100: color_data = 12'b110011110111;
		11'b01101000101: color_data = 12'b110011110111;
		11'b01101000110: color_data = 12'b110011110111;
		11'b01101000111: color_data = 12'b110011110111;
		11'b01101001101: color_data = 12'b110011110111;
		11'b01101001110: color_data = 12'b110011110111;
		11'b01101001111: color_data = 12'b110011110111;
		11'b01101100011: color_data = 12'b110011110111;
		11'b01101100100: color_data = 12'b110011110111;
		11'b01110000100: color_data = 12'b110011110111;
		11'b01110000101: color_data = 12'b110011110111;
		11'b01110000110: color_data = 12'b110011110111;
		11'b01110000111: color_data = 12'b110011110111;
		11'b01110001101: color_data = 12'b110011110111;
		11'b01110001110: color_data = 12'b110011110111;
		11'b01110001111: color_data = 12'b110011110111;
		11'b01110011001: color_data = 12'b110011110111;
		11'b01110100011: color_data = 12'b110011110111;
		11'b01110100100: color_data = 12'b110011110111;
		11'b01111000100: color_data = 12'b110011110111;
		11'b01111000101: color_data = 12'b110011110111;
		11'b01111000110: color_data = 12'b110011110111;
		11'b01111000111: color_data = 12'b110011110111;
		11'b01111001101: color_data = 12'b110011110111;
		11'b01111001110: color_data = 12'b110011110111;
		11'b01111001111: color_data = 12'b110011110111;
		11'b01111010110: color_data = 12'b110011110111;
		11'b01111010111: color_data = 12'b110011110111;
		11'b01111011001: color_data = 12'b110011110111;
		11'b01111011010: color_data = 12'b110011110111;
		11'b01111100010: color_data = 12'b110011110111;
		11'b01111100011: color_data = 12'b110011110111;
		11'b01111100100: color_data = 12'b110011110111;
		11'b10000000100: color_data = 12'b110011110111;
		11'b10000000101: color_data = 12'b110011110111;
		11'b10000000110: color_data = 12'b110011110111;
		11'b10000000111: color_data = 12'b110011110111;
		11'b10000001101: color_data = 12'b110011110111;
		11'b10000001110: color_data = 12'b110011110111;
		11'b10000001111: color_data = 12'b110011110111;
		11'b10000010000: color_data = 12'b110011110111;
		11'b10000010001: color_data = 12'b110011110111;
		11'b10000010010: color_data = 12'b110011110111;
		11'b10000010011: color_data = 12'b110011110111;
		11'b10000010100: color_data = 12'b110011110111;
		11'b10000010101: color_data = 12'b110011110111;
		11'b10000010110: color_data = 12'b110011110111;
		11'b10000011010: color_data = 12'b110011110111;
		11'b10000011011: color_data = 12'b110011110111;
		11'b10000011100: color_data = 12'b110011110111;
		11'b10000011101: color_data = 12'b110011110111;
		11'b10000011110: color_data = 12'b110011110111;
		11'b10000011111: color_data = 12'b110011110111;
		11'b10000100000: color_data = 12'b110011110111;
		11'b10000100001: color_data = 12'b110011110111;
		11'b10000100010: color_data = 12'b110011110111;
		11'b10001000100: color_data = 12'b110011110111;
		11'b10001000101: color_data = 12'b110011110111;
		11'b10001000110: color_data = 12'b110011110111;
		11'b10001000111: color_data = 12'b110011110111;
		11'b10001001101: color_data = 12'b110011110111;
		11'b10001001110: color_data = 12'b110011110111;
		11'b10001001111: color_data = 12'b110011110111;
		11'b10001010000: color_data = 12'b110011110111;
		11'b10001010001: color_data = 12'b110011110111;
		11'b10001010010: color_data = 12'b110011110111;
		11'b10001010011: color_data = 12'b110011110111;
		11'b10001010100: color_data = 12'b110011110111;
		11'b10001010101: color_data = 12'b110011110111;
		11'b10001010110: color_data = 12'b110011110111;
		11'b10001011011: color_data = 12'b110011110111;
		11'b10001011100: color_data = 12'b110011110111;
		11'b10001011101: color_data = 12'b110011110111;
		11'b10001011110: color_data = 12'b110011110111;
		11'b10001011111: color_data = 12'b110011110111;
		11'b10001100000: color_data = 12'b110011110111;
		11'b10001100001: color_data = 12'b110011110111;
		default: color_data = 12'b000000000000;
	endcase
endmodule