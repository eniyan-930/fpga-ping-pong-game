`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.01.2025 14:38:02
// Design Name: 
// Module Name: score_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module score_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		11'b00000000000: color_data = 12'b001110100111;
		11'b00000000001: color_data = 12'b001110100111;
		11'b00000000010: color_data = 12'b001110100111;
		11'b00000000011: color_data = 12'b001110100111;
		11'b00000000100: color_data = 12'b001110100111;
		11'b00000000101: color_data = 12'b001110100111;
		11'b00000000110: color_data = 12'b001110100111;
		11'b00000000111: color_data = 12'b001110100111;
		11'b00000001000: color_data = 12'b001110100111;
		11'b00000001010: color_data = 12'b001110100111;
		11'b00000001011: color_data = 12'b001110100111;
		11'b00000001100: color_data = 12'b001110100111;
		11'b00000001101: color_data = 12'b001110100111;
		11'b00000001110: color_data = 12'b001110100111;
		11'b00000001111: color_data = 12'b001110100111;
		11'b00000010000: color_data = 12'b001110100111;
		11'b00000010001: color_data = 12'b001110100111;
		11'b00000010100: color_data = 12'b001110100111;
		11'b00000010101: color_data = 12'b001110100111;
		11'b00000010110: color_data = 12'b001110100111;
		11'b00000010111: color_data = 12'b001110100111;
		11'b00000011000: color_data = 12'b001110100111;
		11'b00000011001: color_data = 12'b001110100111;
		11'b00000011010: color_data = 12'b001110100111;
		11'b00000011011: color_data = 12'b001110100111;
		11'b00000011110: color_data = 12'b001110100111;
		11'b00000011111: color_data = 12'b001110100111;
		11'b00000100000: color_data = 12'b001110100111;
		11'b00000100001: color_data = 12'b001110100111;
		11'b00000100010: color_data = 12'b001110100111;
		11'b00000100011: color_data = 12'b001110100111;
		11'b00000100100: color_data = 12'b001110100111;
		11'b00000100101: color_data = 12'b001110100111;
		11'b00000101000: color_data = 12'b001110100111;
		11'b00000101001: color_data = 12'b001110100111;
		11'b00000101010: color_data = 12'b001110100111;
		11'b00000101011: color_data = 12'b001110100111;
		11'b00000101100: color_data = 12'b001110100111;
		11'b00000101101: color_data = 12'b001110100111;
		11'b00000101110: color_data = 12'b001110100111;
		11'b00000101111: color_data = 12'b001110100111;
		11'b00001000000: color_data = 12'b001110100111;
		11'b00001000001: color_data = 12'b001110100111;
		11'b00001000010: color_data = 12'b001110100111;
		11'b00001000011: color_data = 12'b001110100111;
		11'b00001000100: color_data = 12'b001110100111;
		11'b00001000101: color_data = 12'b001110100111;
		11'b00001000110: color_data = 12'b001110100111;
		11'b00001000111: color_data = 12'b001110100111;
		11'b00001001000: color_data = 12'b001110100111;
		11'b00001001010: color_data = 12'b001110100111;
		11'b00001001011: color_data = 12'b001110100111;
		11'b00001001100: color_data = 12'b001110100111;
		11'b00001001101: color_data = 12'b001110100111;
		11'b00001001110: color_data = 12'b001110100111;
		11'b00001001111: color_data = 12'b001110100111;
		11'b00001010000: color_data = 12'b001110100111;
		11'b00001010001: color_data = 12'b001110100111;
		11'b00001010100: color_data = 12'b001110100111;
		11'b00001010101: color_data = 12'b001110100111;
		11'b00001010110: color_data = 12'b001110100111;
		11'b00001010111: color_data = 12'b001110100111;
		11'b00001011000: color_data = 12'b001110100111;
		11'b00001011001: color_data = 12'b001110100111;
		11'b00001011010: color_data = 12'b001110100111;
		11'b00001011011: color_data = 12'b001110100111;
		11'b00001011110: color_data = 12'b001110100111;
		11'b00001011111: color_data = 12'b001110100111;
		11'b00001100000: color_data = 12'b001110100111;
		11'b00001100001: color_data = 12'b001110100111;
		11'b00001100010: color_data = 12'b001110100111;
		11'b00001100011: color_data = 12'b001110100111;
		11'b00001100100: color_data = 12'b001110100111;
		11'b00001100101: color_data = 12'b001110100111;
		11'b00001101000: color_data = 12'b001110100111;
		11'b00001101001: color_data = 12'b001110100111;
		11'b00001101010: color_data = 12'b001110100111;
		11'b00001101011: color_data = 12'b001110100111;
		11'b00001101100: color_data = 12'b001110100111;
		11'b00001101101: color_data = 12'b001110100111;
		11'b00001101110: color_data = 12'b001110100111;
		11'b00001101111: color_data = 12'b001110100111;
		11'b00010000000: color_data = 12'b001110100111;
		11'b00010000001: color_data = 12'b001110100111;
		11'b00010000010: color_data = 12'b001110100111;
		11'b00010000011: color_data = 12'b001110100111;
		11'b00010000100: color_data = 12'b001110100111;
		11'b00010000101: color_data = 12'b001110100111;
		11'b00010000110: color_data = 12'b001110100111;
		11'b00010000111: color_data = 12'b001110100111;
		11'b00010001000: color_data = 12'b001110100111;
		11'b00010001010: color_data = 12'b001110100111;
		11'b00010001011: color_data = 12'b001110100111;
		11'b00010001100: color_data = 12'b001110100111;
		11'b00010001101: color_data = 12'b001110100111;
		11'b00010001110: color_data = 12'b001110100111;
		11'b00010001111: color_data = 12'b001110100111;
		11'b00010010000: color_data = 12'b001110100111;
		11'b00010010001: color_data = 12'b001110100111;
		11'b00010010100: color_data = 12'b001110100111;
		11'b00010010101: color_data = 12'b001110100111;
		11'b00010010110: color_data = 12'b001110100111;
		11'b00010010111: color_data = 12'b001110100111;
		11'b00010011000: color_data = 12'b001110100111;
		11'b00010011001: color_data = 12'b001110100111;
		11'b00010011010: color_data = 12'b001110100111;
		11'b00010011011: color_data = 12'b001110100111;
		11'b00010011110: color_data = 12'b001110100111;
		11'b00010011111: color_data = 12'b001110100111;
		11'b00010100000: color_data = 12'b001110100111;
		11'b00010100001: color_data = 12'b001110100111;
		11'b00010100010: color_data = 12'b001110100111;
		11'b00010100011: color_data = 12'b001110100111;
		11'b00010100100: color_data = 12'b001110100111;
		11'b00010100101: color_data = 12'b001110100111;
		11'b00010101000: color_data = 12'b001110100111;
		11'b00010101001: color_data = 12'b001110100111;
		11'b00010101010: color_data = 12'b001110100111;
		11'b00010101011: color_data = 12'b001110100111;
		11'b00010101100: color_data = 12'b001110100111;
		11'b00010101101: color_data = 12'b001110100111;
		11'b00010101110: color_data = 12'b001110100111;
		11'b00010101111: color_data = 12'b001110100111;
		11'b00011000000: color_data = 12'b001110100111;
		11'b00011000001: color_data = 12'b001110100111;
		11'b00011000010: color_data = 12'b001110100111;
		11'b00011001010: color_data = 12'b001110100111;
		11'b00011001011: color_data = 12'b001110100111;
		11'b00011010100: color_data = 12'b001110100111;
		11'b00011010101: color_data = 12'b001110100111;
		11'b00011011010: color_data = 12'b001110100111;
		11'b00011011011: color_data = 12'b001110100111;
		11'b00011011110: color_data = 12'b001110100111;
		11'b00011011111: color_data = 12'b001110100111;
		11'b00011100100: color_data = 12'b001110100111;
		11'b00011100101: color_data = 12'b001110100111;
		11'b00011101000: color_data = 12'b001110100111;
		11'b00011101001: color_data = 12'b001110100111;
		11'b00100000000: color_data = 12'b001110100111;
		11'b00100000001: color_data = 12'b001110100111;
		11'b00100000010: color_data = 12'b001110100111;
		11'b00100001010: color_data = 12'b001110100111;
		11'b00100001011: color_data = 12'b001110100111;
		11'b00100010100: color_data = 12'b001110100111;
		11'b00100010101: color_data = 12'b001110100111;
		11'b00100011010: color_data = 12'b001110100111;
		11'b00100011011: color_data = 12'b001110100111;
		11'b00100011110: color_data = 12'b001110100111;
		11'b00100011111: color_data = 12'b001110100111;
		11'b00100100100: color_data = 12'b001110100111;
		11'b00100100101: color_data = 12'b001110100111;
		11'b00100101000: color_data = 12'b001110100111;
		11'b00100101001: color_data = 12'b001110100111;
		11'b00101000000: color_data = 12'b001110100111;
		11'b00101000001: color_data = 12'b001110100111;
		11'b00101000010: color_data = 12'b001110100111;
		11'b00101001010: color_data = 12'b001110100111;
		11'b00101001011: color_data = 12'b001110100111;
		11'b00101010100: color_data = 12'b001110100111;
		11'b00101010101: color_data = 12'b001110100111;
		11'b00101011010: color_data = 12'b001110100111;
		11'b00101011011: color_data = 12'b001110100111;
		11'b00101011110: color_data = 12'b001110100111;
		11'b00101011111: color_data = 12'b001110100111;
		11'b00101100100: color_data = 12'b001110100111;
		11'b00101100101: color_data = 12'b001110100111;
		11'b00101101000: color_data = 12'b001110100111;
		11'b00101101001: color_data = 12'b001110100111;
		11'b00101110101: color_data = 12'b001110100111;
		11'b00101110110: color_data = 12'b001110100111;
		11'b00101110111: color_data = 12'b001110100111;
		11'b00110000000: color_data = 12'b001110100111;
		11'b00110000001: color_data = 12'b001110100111;
		11'b00110000010: color_data = 12'b001110100111;
		11'b00110001010: color_data = 12'b001110100111;
		11'b00110001011: color_data = 12'b001110100111;
		11'b00110010100: color_data = 12'b001110100111;
		11'b00110010101: color_data = 12'b001110100111;
		11'b00110011010: color_data = 12'b001110100111;
		11'b00110011011: color_data = 12'b001110100111;
		11'b00110011110: color_data = 12'b001110100111;
		11'b00110011111: color_data = 12'b001110100111;
		11'b00110100100: color_data = 12'b001110100111;
		11'b00110100101: color_data = 12'b001110100111;
		11'b00110101000: color_data = 12'b001110100111;
		11'b00110101001: color_data = 12'b001110100111;
		11'b00110110101: color_data = 12'b001110100111;
		11'b00110110110: color_data = 12'b001110100111;
		11'b00110110111: color_data = 12'b001110100111;
		11'b00111000000: color_data = 12'b001110100111;
		11'b00111000001: color_data = 12'b001110100111;
		11'b00111000010: color_data = 12'b001110100111;
		11'b00111000011: color_data = 12'b001110100111;
		11'b00111000100: color_data = 12'b001110100111;
		11'b00111000101: color_data = 12'b001110100111;
		11'b00111000110: color_data = 12'b001110100111;
		11'b00111000111: color_data = 12'b001110100111;
		11'b00111001000: color_data = 12'b001110100111;
		11'b00111001010: color_data = 12'b001110100111;
		11'b00111001011: color_data = 12'b001110100111;
		11'b00111010100: color_data = 12'b001110100111;
		11'b00111010101: color_data = 12'b001110100111;
		11'b00111011010: color_data = 12'b001110100111;
		11'b00111011011: color_data = 12'b001110100111;
		11'b00111011110: color_data = 12'b001110100111;
		11'b00111011111: color_data = 12'b001110100111;
		11'b00111100000: color_data = 12'b001110100111;
		11'b00111100001: color_data = 12'b001110100111;
		11'b00111100010: color_data = 12'b001110100111;
		11'b00111100011: color_data = 12'b001110100111;
		11'b00111101000: color_data = 12'b001110100111;
		11'b00111101001: color_data = 12'b001110100111;
		11'b00111101010: color_data = 12'b001110100111;
		11'b00111101011: color_data = 12'b001110100111;
		11'b00111101100: color_data = 12'b001110100111;
		11'b00111101101: color_data = 12'b001110100111;
		11'b00111101110: color_data = 12'b001110100111;
		11'b00111101111: color_data = 12'b001110100111;
		11'b00111110101: color_data = 12'b001110100111;
		11'b00111110110: color_data = 12'b001110100111;
		11'b00111110111: color_data = 12'b001110100111;
		11'b01000000000: color_data = 12'b001110100111;
		11'b01000000001: color_data = 12'b001110100111;
		11'b01000000010: color_data = 12'b001110100111;
		11'b01000000011: color_data = 12'b001110100111;
		11'b01000000100: color_data = 12'b001110100111;
		11'b01000000101: color_data = 12'b001110100111;
		11'b01000000110: color_data = 12'b001110100111;
		11'b01000000111: color_data = 12'b001110100111;
		11'b01000001000: color_data = 12'b001110100111;
		11'b01000001010: color_data = 12'b001110100111;
		11'b01000001011: color_data = 12'b001110100111;
		11'b01000010100: color_data = 12'b001110100111;
		11'b01000010101: color_data = 12'b001110100111;
		11'b01000011010: color_data = 12'b001110100111;
		11'b01000011011: color_data = 12'b001110100111;
		11'b01000011110: color_data = 12'b001110100111;
		11'b01000011111: color_data = 12'b001110100111;
		11'b01000100000: color_data = 12'b001110100111;
		11'b01000100001: color_data = 12'b001110100111;
		11'b01000100010: color_data = 12'b001110100111;
		11'b01000100011: color_data = 12'b001110100111;
		11'b01000101000: color_data = 12'b001110100111;
		11'b01000101001: color_data = 12'b001110100111;
		11'b01000101010: color_data = 12'b001110100111;
		11'b01000101011: color_data = 12'b001110100111;
		11'b01000101100: color_data = 12'b001110100111;
		11'b01000101101: color_data = 12'b001110100111;
		11'b01000101110: color_data = 12'b001110100111;
		11'b01000101111: color_data = 12'b001110100111;
		11'b01001000000: color_data = 12'b001110100111;
		11'b01001000001: color_data = 12'b001110100111;
		11'b01001000010: color_data = 12'b001110100111;
		11'b01001000011: color_data = 12'b001110100111;
		11'b01001000100: color_data = 12'b001110100111;
		11'b01001000101: color_data = 12'b001110100111;
		11'b01001000110: color_data = 12'b001110100111;
		11'b01001000111: color_data = 12'b001110100111;
		11'b01001001000: color_data = 12'b001110100111;
		11'b01001001010: color_data = 12'b001110100111;
		11'b01001001011: color_data = 12'b001110100111;
		11'b01001010100: color_data = 12'b001110100111;
		11'b01001010101: color_data = 12'b001110100111;
		11'b01001011010: color_data = 12'b001110100111;
		11'b01001011011: color_data = 12'b001110100111;
		11'b01001011110: color_data = 12'b001110100111;
		11'b01001011111: color_data = 12'b001110100111;
		11'b01001100000: color_data = 12'b001110100111;
		11'b01001100001: color_data = 12'b001110100111;
		11'b01001100010: color_data = 12'b001110100111;
		11'b01001100011: color_data = 12'b001110100111;
		11'b01001101000: color_data = 12'b001110100111;
		11'b01001101001: color_data = 12'b001110100111;
		11'b01001101010: color_data = 12'b001110100111;
		11'b01001101011: color_data = 12'b001110100111;
		11'b01001101100: color_data = 12'b001110100111;
		11'b01001101101: color_data = 12'b001110100111;
		11'b01001101110: color_data = 12'b001110100111;
		11'b01001101111: color_data = 12'b001110100111;
		11'b01010000000: color_data = 12'b001110100111;
		11'b01010000001: color_data = 12'b001110100111;
		11'b01010000010: color_data = 12'b001110100111;
		11'b01010000011: color_data = 12'b001110100111;
		11'b01010000100: color_data = 12'b001110100111;
		11'b01010000101: color_data = 12'b001110100111;
		11'b01010000110: color_data = 12'b001110100111;
		11'b01010000111: color_data = 12'b001110100111;
		11'b01010001000: color_data = 12'b001110100111;
		11'b01010001010: color_data = 12'b001110100111;
		11'b01010001011: color_data = 12'b001110100111;
		11'b01010010100: color_data = 12'b001110100111;
		11'b01010010101: color_data = 12'b001110100111;
		11'b01010011010: color_data = 12'b001110100111;
		11'b01010011011: color_data = 12'b001110100111;
		11'b01010011110: color_data = 12'b001110100111;
		11'b01010011111: color_data = 12'b001110100111;
		11'b01010100000: color_data = 12'b001110100111;
		11'b01010100001: color_data = 12'b001110100111;
		11'b01010100010: color_data = 12'b001110100111;
		11'b01010100011: color_data = 12'b001110100111;
		11'b01010101000: color_data = 12'b001110100111;
		11'b01010101001: color_data = 12'b001110100111;
		11'b01010101010: color_data = 12'b001110100111;
		11'b01010101011: color_data = 12'b001110100111;
		11'b01010101100: color_data = 12'b001110100111;
		11'b01010101101: color_data = 12'b001110100111;
		11'b01010101110: color_data = 12'b001110100111;
		11'b01010101111: color_data = 12'b001110100111;
		11'b01011000110: color_data = 12'b001110100111;
		11'b01011000111: color_data = 12'b001110100111;
		11'b01011001000: color_data = 12'b001110100111;
		11'b01011001010: color_data = 12'b001110100111;
		11'b01011001011: color_data = 12'b001110100111;
		11'b01011010100: color_data = 12'b001110100111;
		11'b01011010101: color_data = 12'b001110100111;
		11'b01011011010: color_data = 12'b001110100111;
		11'b01011011011: color_data = 12'b001110100111;
		11'b01011011110: color_data = 12'b001110100111;
		11'b01011011111: color_data = 12'b001110100111;
		11'b01011100100: color_data = 12'b001110100111;
		11'b01011100101: color_data = 12'b001110100111;
		11'b01011101000: color_data = 12'b001110100111;
		11'b01011101001: color_data = 12'b001110100111;
		11'b01011110101: color_data = 12'b001110100111;
		11'b01011110110: color_data = 12'b001110100111;
		11'b01011110111: color_data = 12'b001110100111;
		11'b01100000110: color_data = 12'b001110100111;
		11'b01100000111: color_data = 12'b001110100111;
		11'b01100001000: color_data = 12'b001110100111;
		11'b01100001010: color_data = 12'b001110100111;
		11'b01100001011: color_data = 12'b001110100111;
		11'b01100010100: color_data = 12'b001110100111;
		11'b01100010101: color_data = 12'b001110100111;
		11'b01100011010: color_data = 12'b001110100111;
		11'b01100011011: color_data = 12'b001110100111;
		11'b01100011110: color_data = 12'b001110100111;
		11'b01100011111: color_data = 12'b001110100111;
		11'b01100100100: color_data = 12'b001110100111;
		11'b01100100101: color_data = 12'b001110100111;
		11'b01100101000: color_data = 12'b001110100111;
		11'b01100101001: color_data = 12'b001110100111;
		11'b01100110101: color_data = 12'b001110100111;
		11'b01100110110: color_data = 12'b001110100111;
		11'b01100110111: color_data = 12'b001110100111;
		11'b01101000110: color_data = 12'b001110100111;
		11'b01101000111: color_data = 12'b001110100111;
		11'b01101001000: color_data = 12'b001110100111;
		11'b01101001010: color_data = 12'b001110100111;
		11'b01101001011: color_data = 12'b001110100111;
		11'b01101010100: color_data = 12'b001110100111;
		11'b01101010101: color_data = 12'b001110100111;
		11'b01101011010: color_data = 12'b001110100111;
		11'b01101011011: color_data = 12'b001110100111;
		11'b01101011110: color_data = 12'b001110100111;
		11'b01101011111: color_data = 12'b001110100111;
		11'b01101100100: color_data = 12'b001110100111;
		11'b01101100101: color_data = 12'b001110100111;
		11'b01101101000: color_data = 12'b001110100111;
		11'b01101101001: color_data = 12'b001110100111;
		11'b01101110101: color_data = 12'b001110100111;
		11'b01101110110: color_data = 12'b001110100111;
		11'b01101110111: color_data = 12'b001110100111;
		11'b01110000110: color_data = 12'b001110100111;
		11'b01110000111: color_data = 12'b001110100111;
		11'b01110001000: color_data = 12'b001110100111;
		11'b01110001010: color_data = 12'b001110100111;
		11'b01110001011: color_data = 12'b001110100111;
		11'b01110010100: color_data = 12'b001110100111;
		11'b01110010101: color_data = 12'b001110100111;
		11'b01110011010: color_data = 12'b001110100111;
		11'b01110011011: color_data = 12'b001110100111;
		11'b01110011110: color_data = 12'b001110100111;
		11'b01110011111: color_data = 12'b001110100111;
		11'b01110100100: color_data = 12'b001110100111;
		11'b01110100101: color_data = 12'b001110100111;
		11'b01110101000: color_data = 12'b001110100111;
		11'b01110101001: color_data = 12'b001110100111;
		11'b01111000000: color_data = 12'b001110100111;
		11'b01111000001: color_data = 12'b001110100111;
		11'b01111000010: color_data = 12'b001110100111;
		11'b01111000011: color_data = 12'b001110100111;
		11'b01111000100: color_data = 12'b001110100111;
		11'b01111000101: color_data = 12'b001110100111;
		11'b01111000110: color_data = 12'b001110100111;
		11'b01111000111: color_data = 12'b001110100111;
		11'b01111001000: color_data = 12'b001110100111;
		11'b01111001010: color_data = 12'b001110100111;
		11'b01111001011: color_data = 12'b001110100111;
		11'b01111001100: color_data = 12'b001110100111;
		11'b01111001101: color_data = 12'b001110100111;
		11'b01111001110: color_data = 12'b001110100111;
		11'b01111001111: color_data = 12'b001110100111;
		11'b01111010000: color_data = 12'b001110100111;
		11'b01111010001: color_data = 12'b001110100111;
		11'b01111010100: color_data = 12'b001110100111;
		11'b01111010101: color_data = 12'b001110100111;
		11'b01111010110: color_data = 12'b001110100111;
		11'b01111010111: color_data = 12'b001110100111;
		11'b01111011000: color_data = 12'b001110100111;
		11'b01111011001: color_data = 12'b001110100111;
		11'b01111011010: color_data = 12'b001110100111;
		11'b01111011011: color_data = 12'b001110100111;
		11'b01111011110: color_data = 12'b001110100111;
		11'b01111011111: color_data = 12'b001110100111;
		11'b01111100100: color_data = 12'b001110100111;
		11'b01111100101: color_data = 12'b001110100111;
		11'b01111101000: color_data = 12'b001110100111;
		11'b01111101001: color_data = 12'b001110100111;
		11'b01111101010: color_data = 12'b001110100111;
		11'b01111101011: color_data = 12'b001110100111;
		11'b01111101100: color_data = 12'b001110100111;
		11'b01111101101: color_data = 12'b001110100111;
		11'b01111101110: color_data = 12'b001110100111;
		11'b01111101111: color_data = 12'b001110100111;
		11'b10000000000: color_data = 12'b001110100111;
		11'b10000000001: color_data = 12'b001110100111;
		11'b10000000010: color_data = 12'b001110100111;
		11'b10000000011: color_data = 12'b001110100111;
		11'b10000000100: color_data = 12'b001110100111;
		11'b10000000101: color_data = 12'b001110100111;
		11'b10000000110: color_data = 12'b001110100111;
		11'b10000000111: color_data = 12'b001110100111;
		11'b10000001000: color_data = 12'b001110100111;
		11'b10000001010: color_data = 12'b001110100111;
		11'b10000001011: color_data = 12'b001110100111;
		11'b10000001100: color_data = 12'b001110100111;
		11'b10000001101: color_data = 12'b001110100111;
		11'b10000001110: color_data = 12'b001110100111;
		11'b10000001111: color_data = 12'b001110100111;
		11'b10000010000: color_data = 12'b001110100111;
		11'b10000010001: color_data = 12'b001110100111;
		11'b10000010100: color_data = 12'b001110100111;
		11'b10000010101: color_data = 12'b001110100111;
		11'b10000010110: color_data = 12'b001110100111;
		11'b10000010111: color_data = 12'b001110100111;
		11'b10000011000: color_data = 12'b001110100111;
		11'b10000011001: color_data = 12'b001110100111;
		11'b10000011010: color_data = 12'b001110100111;
		11'b10000011011: color_data = 12'b001110100111;
		11'b10000011110: color_data = 12'b001110100111;
		11'b10000011111: color_data = 12'b001110100111;
		11'b10000100100: color_data = 12'b001110100111;
		11'b10000100101: color_data = 12'b001110100111;
		11'b10000101000: color_data = 12'b001110100111;
		11'b10000101001: color_data = 12'b001110100111;
		11'b10000101010: color_data = 12'b001110100111;
		11'b10000101011: color_data = 12'b001110100111;
		11'b10000101100: color_data = 12'b001110100111;
		11'b10000101101: color_data = 12'b001110100111;
		11'b10000101110: color_data = 12'b001110100111;
		11'b10000101111: color_data = 12'b001110100111;
		11'b10001000000: color_data = 12'b001110100111;
		11'b10001000001: color_data = 12'b001110100111;
		11'b10001000010: color_data = 12'b001110100111;
		11'b10001000011: color_data = 12'b001110100111;
		11'b10001000100: color_data = 12'b001110100111;
		11'b10001000101: color_data = 12'b001110100111;
		11'b10001000110: color_data = 12'b001110100111;
		11'b10001000111: color_data = 12'b001110100111;
		11'b10001001000: color_data = 12'b001110100111;
		11'b10001001010: color_data = 12'b001110100111;
		11'b10001001011: color_data = 12'b001110100111;
		11'b10001001100: color_data = 12'b001110100111;
		11'b10001001101: color_data = 12'b001110100111;
		11'b10001001110: color_data = 12'b001110100111;
		11'b10001001111: color_data = 12'b001110100111;
		11'b10001010000: color_data = 12'b001110100111;
		11'b10001010001: color_data = 12'b001110100111;
		11'b10001010100: color_data = 12'b001110100111;
		11'b10001010101: color_data = 12'b001110100111;
		11'b10001010110: color_data = 12'b001110100111;
		11'b10001010111: color_data = 12'b001110100111;
		11'b10001011000: color_data = 12'b001110100111;
		11'b10001011001: color_data = 12'b001110100111;
		11'b10001011010: color_data = 12'b001110100111;
		11'b10001011011: color_data = 12'b001110100111;
		11'b10001011110: color_data = 12'b001110100111;
		11'b10001011111: color_data = 12'b001110100111;
		11'b10001100100: color_data = 12'b001110100111;
		11'b10001100101: color_data = 12'b001110100111;
		11'b10001101000: color_data = 12'b001110100111;
		11'b10001101001: color_data = 12'b001110100111;
		11'b10001101010: color_data = 12'b001110100111;
		11'b10001101011: color_data = 12'b001110100111;
		11'b10001101100: color_data = 12'b001110100111;
		11'b10001101101: color_data = 12'b001110100111;
		11'b10001101110: color_data = 12'b001110100111;
		11'b10001101111: color_data = 12'b001110100111;
		default: color_data  = 12'b000000000000;
	endcase
endmodule
