`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.01.2025 14:36:52
// Design Name: 
// Module Name: number_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module number_rom
	(
		input wire clk,
		input wire [3:0] row,
		input wire [3:0] col,
        input wire [3:0] score,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [3:0] row_reg;
	reg [3:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({score,row_reg, col_reg})
		12'b000000000011: color_data = 12'b001110100111;
		12'b000000000100: color_data = 12'b001110100111;
		12'b000000000101: color_data = 12'b001110100111;
		12'b000000000110: color_data = 12'b001110100111;
		12'b000000000111: color_data = 12'b001110100111;
		12'b000000001000: color_data = 12'b001110100111;
		12'b000000001001: color_data = 12'b001110100111;
		12'b000000001010: color_data = 12'b001110100111;
		12'b000000010011: color_data = 12'b001110100111;
		12'b000000010100: color_data = 12'b001110100111;
		12'b000000010101: color_data = 12'b001110100111;
		12'b000000010110: color_data = 12'b001110100111;
		12'b000000010111: color_data = 12'b001110100111;
		12'b000000011000: color_data = 12'b001110100111;
		12'b000000011001: color_data = 12'b001110100111;
		12'b000000011010: color_data = 12'b001110100111;
		12'b000000100000: color_data = 12'b001110100111;
		12'b000000100001: color_data = 12'b001110100111;
		12'b000000100010: color_data = 12'b001110100111;
		12'b000000101011: color_data = 12'b001110100111;
		12'b000000101100: color_data = 12'b001110100111;
		12'b000000110000: color_data = 12'b001110100111;
		12'b000000110001: color_data = 12'b001110100111;
		12'b000000110010: color_data = 12'b001110100111;
		12'b000000111011: color_data = 12'b001110100111;
		12'b000000111100: color_data = 12'b001110100111;
		12'b000001000000: color_data = 12'b001110100111;
		12'b000001000001: color_data = 12'b001110100111;
		12'b000001000010: color_data = 12'b001110100111;
		12'b000001001011: color_data = 12'b001110100111;
		12'b000001001100: color_data = 12'b001110100111;
		12'b000001010000: color_data = 12'b001110100111;
		12'b000001010001: color_data = 12'b001110100111;
		12'b000001010010: color_data = 12'b001110100111;
		12'b000001011011: color_data = 12'b001110100111;
		12'b000001011100: color_data = 12'b001110100111;
		12'b000001100000: color_data = 12'b001110100111;
		12'b000001100001: color_data = 12'b001110100111;
		12'b000001100010: color_data = 12'b001110100111;
		12'b000001101011: color_data = 12'b001110100111;
		12'b000001101100: color_data = 12'b001110100111;
		12'b000001110000: color_data = 12'b001110100111;
		12'b000001110001: color_data = 12'b001110100111;
		12'b000001110010: color_data = 12'b001110100111;
		12'b000001111011: color_data = 12'b001110100111;
		12'b000001111100: color_data = 12'b001110100111;
		12'b000010000000: color_data = 12'b001110100111;
		12'b000010000001: color_data = 12'b001110100111;
		12'b000010000010: color_data = 12'b001110100111;
		12'b000010001011: color_data = 12'b001110100111;
		12'b000010001100: color_data = 12'b001110100111;
		12'b000010010000: color_data = 12'b001110100111;
		12'b000010010001: color_data = 12'b001110100111;
		12'b000010010010: color_data = 12'b001110100111;
		12'b000010011011: color_data = 12'b001110100111;
		12'b000010011100: color_data = 12'b001110100111;
		12'b000010100000: color_data = 12'b001110100111;
		12'b000010100001: color_data = 12'b001110100111;
		12'b000010100010: color_data = 12'b001110100111;
		12'b000010101011: color_data = 12'b001110100111;
		12'b000010101100: color_data = 12'b001110100111;
		12'b000010110000: color_data = 12'b001110100111;
		12'b000010110001: color_data = 12'b001110100111;
		12'b000010110010: color_data = 12'b001110100111;
		12'b000010111011: color_data = 12'b001110100111;
		12'b000010111100: color_data = 12'b001110100111;
		12'b000011000011: color_data = 12'b001110100111;
		12'b000011000100: color_data = 12'b001110100111;
		12'b000011000101: color_data = 12'b001110100111;
		12'b000011000110: color_data = 12'b001110100111;
		12'b000011000111: color_data = 12'b001110100111;
		12'b000011001000: color_data = 12'b001110100111;
		12'b000011001001: color_data = 12'b001110100111;
		12'b000011001010: color_data = 12'b001110100111;
		12'b000011010011: color_data = 12'b001110100111;
		12'b000011010100: color_data = 12'b001110100111;
		12'b000011010101: color_data = 12'b001110100111;
		12'b000011010110: color_data = 12'b001110100111;
		12'b000011010111: color_data = 12'b001110100111;
		12'b000011011000: color_data = 12'b001110100111;
		12'b000011011001: color_data = 12'b001110100111;
		12'b000011011010: color_data = 12'b001110100111;
        12'b000100000110: color_data = 12'b001110100111;
		12'b000100000111: color_data = 12'b001110100111;
		12'b000100010110: color_data = 12'b001110100111;
		12'b000100010111: color_data = 12'b001110100111;
		12'b000100100011: color_data = 12'b001110100111;
		12'b000100100100: color_data = 12'b001110100111;
		12'b000100100101: color_data = 12'b001110100111;
		12'b000100100110: color_data = 12'b001110100111;
		12'b000100100111: color_data = 12'b001110100111;
		12'b000100110011: color_data = 12'b001110100111;
		12'b000100110100: color_data = 12'b001110100111;
		12'b000100110101: color_data = 12'b001110100111;
		12'b000100110110: color_data = 12'b001110100111;
		12'b000100110111: color_data = 12'b001110100111;
		12'b000101000110: color_data = 12'b001110100111;
		12'b000101000111: color_data = 12'b001110100111;
		12'b000101010110: color_data = 12'b001110100111;
		12'b000101010111: color_data = 12'b001110100111;
		12'b000101100110: color_data = 12'b001110100111;
		12'b000101100111: color_data = 12'b001110100111;
		12'b000101110110: color_data = 12'b001110100111;
		12'b000101110111: color_data = 12'b001110100111;
		12'b000110000110: color_data = 12'b001110100111;
		12'b000110000111: color_data = 12'b001110100111;
		12'b000110010110: color_data = 12'b001110100111;
		12'b000110010111: color_data = 12'b001110100111;
		12'b000110100110: color_data = 12'b001110100111;
		12'b000110100111: color_data = 12'b001110100111;
		12'b000110110110: color_data = 12'b001110100111;
		12'b000110110111: color_data = 12'b001110100111;
		12'b000111000000: color_data = 12'b001110100111;
		12'b000111000001: color_data = 12'b001110100111;
		12'b000111000010: color_data = 12'b001110100111;
		12'b000111000011: color_data = 12'b001110100111;
		12'b000111000100: color_data = 12'b001110100111;
		12'b000111000101: color_data = 12'b001110100111;
		12'b000111000110: color_data = 12'b001110100111;
		12'b000111000111: color_data = 12'b001110100111;
		12'b000111001000: color_data = 12'b001110100111;
		12'b000111001001: color_data = 12'b001110100111;
		12'b000111001010: color_data = 12'b001110100111;
		12'b000111001011: color_data = 12'b001110100111;
		12'b000111001100: color_data = 12'b001110100111;
		12'b000111010000: color_data = 12'b001110100111;
		12'b000111010001: color_data = 12'b001110100111;
		12'b000111010010: color_data = 12'b001110100111;
		12'b000111010011: color_data = 12'b001110100111;
		12'b000111010100: color_data = 12'b001110100111;
		12'b000111010101: color_data = 12'b001110100111;
		12'b000111010110: color_data = 12'b001110100111;
		12'b000111010111: color_data = 12'b001110100111;
		12'b000111011000: color_data = 12'b001110100111;
		12'b000111011001: color_data = 12'b001110100111;
		12'b000111011010: color_data = 12'b001110100111;
		12'b000111011011: color_data = 12'b001110100111;
		12'b000111011100: color_data = 12'b001110100111;
        12'b001000000100: color_data = 12'b001110100111;
		12'b001000000101: color_data = 12'b001110100111;
		12'b001000000110: color_data = 12'b001110100111;
		12'b001000000111: color_data = 12'b001110100111;
		12'b001000001000: color_data = 12'b001110100111;
		12'b001000001001: color_data = 12'b001110100111;
		12'b001000001010: color_data = 12'b001110100111;
		12'b001000001011: color_data = 12'b001110100111;
		12'b001000010100: color_data = 12'b001110100111;
		12'b001000010101: color_data = 12'b001110100111;
		12'b001000010110: color_data = 12'b001110100111;
		12'b001000010111: color_data = 12'b001110100111;
		12'b001000011000: color_data = 12'b001110100111;
		12'b001000011001: color_data = 12'b001110100111;
		12'b001000011010: color_data = 12'b001110100111;
		12'b001000011011: color_data = 12'b001110100111;
		12'b001000100000: color_data = 12'b001110100111;
		12'b001000100001: color_data = 12'b001110100111;
		12'b001000100010: color_data = 12'b001110100111;
		12'b001000100011: color_data = 12'b001110100111;
		12'b001000101100: color_data = 12'b001110100111;
		12'b001000110000: color_data = 12'b001110100111;
		12'b001000110001: color_data = 12'b001110100111;
		12'b001000110010: color_data = 12'b001110100111;
		12'b001000110011: color_data = 12'b001110100111;
		12'b001000111100: color_data = 12'b001110100111;
		12'b001001001100: color_data = 12'b001110100111;
		12'b001001011100: color_data = 12'b001110100111;
		12'b001001101001: color_data = 12'b001110100111;
		12'b001001101010: color_data = 12'b001110100111;
		12'b001001101011: color_data = 12'b001110100111;
		12'b001001111001: color_data = 12'b001110100111;
		12'b001001111010: color_data = 12'b001110100111;
		12'b001001111011: color_data = 12'b001110100111;
		12'b001010000111: color_data = 12'b001110100111;
		12'b001010001000: color_data = 12'b001110100111;
		12'b001010010111: color_data = 12'b001110100111;
		12'b001010011000: color_data = 12'b001110100111;
		12'b001010100100: color_data = 12'b001110100111;
		12'b001010100101: color_data = 12'b001110100111;
		12'b001010100110: color_data = 12'b001110100111;
		12'b001010110100: color_data = 12'b001110100111;
		12'b001010110101: color_data = 12'b001110100111;
		12'b001010110110: color_data = 12'b001110100111;
		12'b001011000000: color_data = 12'b001110100111;
		12'b001011000001: color_data = 12'b001110100111;
		12'b001011000010: color_data = 12'b001110100111;
		12'b001011000011: color_data = 12'b001110100111;
		12'b001011000100: color_data = 12'b001110100111;
		12'b001011000101: color_data = 12'b001110100111;
		12'b001011000110: color_data = 12'b001110100111;
		12'b001011000111: color_data = 12'b001110100111;
		12'b001011001000: color_data = 12'b001110100111;
		12'b001011001001: color_data = 12'b001110100111;
		12'b001011001010: color_data = 12'b001110100111;
		12'b001011001011: color_data = 12'b001110100111;
		12'b001011001100: color_data = 12'b001110100111;
		12'b001011010000: color_data = 12'b001110100111;
		12'b001011010001: color_data = 12'b001110100111;
		12'b001011010010: color_data = 12'b001110100111;
		12'b001011010011: color_data = 12'b001110100111;
		12'b001011010100: color_data = 12'b001110100111;
		12'b001011010101: color_data = 12'b001110100111;
		12'b001011010110: color_data = 12'b001110100111;
		12'b001011010111: color_data = 12'b001110100111;
		12'b001011011000: color_data = 12'b001110100111;
		12'b001011011001: color_data = 12'b001110100111;
		12'b001011011010: color_data = 12'b001110100111;
		12'b001011011011: color_data = 12'b001110100111;
		12'b001011011100: color_data = 12'b001110100111;
        12'b001100000011: color_data = 12'b001110100111;
		12'b001100000100: color_data = 12'b001110100111;
		12'b001100000101: color_data = 12'b001110100111;
		12'b001100000110: color_data = 12'b001110100111;
		12'b001100000111: color_data = 12'b001110100111;
		12'b001100001000: color_data = 12'b001110100111;
		12'b001100001001: color_data = 12'b001110100111;
		12'b001100001010: color_data = 12'b001110100111;
		12'b001100010011: color_data = 12'b001110100111;
		12'b001100010100: color_data = 12'b001110100111;
		12'b001100010101: color_data = 12'b001110100111;
		12'b001100010110: color_data = 12'b001110100111;
		12'b001100010111: color_data = 12'b001110100111;
		12'b001100011000: color_data = 12'b001110100111;
		12'b001100011001: color_data = 12'b001110100111;
		12'b001100011010: color_data = 12'b001110100111;
		12'b001100100000: color_data = 12'b001110100111;
		12'b001100100001: color_data = 12'b001110100111;
		12'b001100100010: color_data = 12'b001110100111;
		12'b001100101011: color_data = 12'b001110100111;
		12'b001100101100: color_data = 12'b001110100111;
		12'b001100110000: color_data = 12'b001110100111;
		12'b001100110001: color_data = 12'b001110100111;
		12'b001100110010: color_data = 12'b001110100111;
		12'b001100111011: color_data = 12'b001110100111;
		12'b001100111100: color_data = 12'b001110100111;
		12'b001101001011: color_data = 12'b001110100111;
		12'b001101001100: color_data = 12'b001110100111;
		12'b001101011011: color_data = 12'b001110100111;
		12'b001101011100: color_data = 12'b001110100111;
		12'b001101100110: color_data = 12'b001110100111;
		12'b001101100111: color_data = 12'b001110100111;
		12'b001101101000: color_data = 12'b001110100111;
		12'b001101101001: color_data = 12'b001110100111;
		12'b001101101010: color_data = 12'b001110100111;
		12'b001101110110: color_data = 12'b001110100111;
		12'b001101110111: color_data = 12'b001110100111;
		12'b001101111000: color_data = 12'b001110100111;
		12'b001101111001: color_data = 12'b001110100111;
		12'b001101111010: color_data = 12'b001110100111;
		12'b001110001011: color_data = 12'b001110100111;
		12'b001110001100: color_data = 12'b001110100111;
		12'b001110011011: color_data = 12'b001110100111;
		12'b001110011100: color_data = 12'b001110100111;
		12'b001110100000: color_data = 12'b001110100111;
		12'b001110100001: color_data = 12'b001110100111;
		12'b001110100010: color_data = 12'b001110100111;
		12'b001110101011: color_data = 12'b001110100111;
		12'b001110101100: color_data = 12'b001110100111;
		12'b001110110000: color_data = 12'b001110100111;
		12'b001110110001: color_data = 12'b001110100111;
		12'b001110110010: color_data = 12'b001110100111;
		12'b001110111011: color_data = 12'b001110100111;
		12'b001110111100: color_data = 12'b001110100111;
		12'b001111000011: color_data = 12'b001110100111;
		12'b001111000100: color_data = 12'b001110100111;
		12'b001111000101: color_data = 12'b001110100111;
		12'b001111000110: color_data = 12'b001110100111;
		12'b001111000111: color_data = 12'b001110100111;
		12'b001111001000: color_data = 12'b001110100111;
		12'b001111001001: color_data = 12'b001110100111;
		12'b001111001010: color_data = 12'b001110100111;
		12'b001111010011: color_data = 12'b001110100111;
		12'b001111010100: color_data = 12'b001110100111;
		12'b001111010101: color_data = 12'b001110100111;
		12'b001111010110: color_data = 12'b001110100111;
		12'b001111010111: color_data = 12'b001110100111;
		12'b001111011000: color_data = 12'b001110100111;
		12'b001111011001: color_data = 12'b001110100111;
		12'b001111011010: color_data = 12'b001110100111;
        12'b010000001000: color_data = 12'b001110100111;
		12'b010000001001: color_data = 12'b001110100111;
		12'b010000001010: color_data = 12'b001110100111;
		12'b010000011000: color_data = 12'b001110100111;
		12'b010000011001: color_data = 12'b001110100111;
		12'b010000011010: color_data = 12'b001110100111;
		12'b010000100110: color_data = 12'b001110100111;
		12'b010000100111: color_data = 12'b001110100111;
		12'b010000101000: color_data = 12'b001110100111;
		12'b010000101001: color_data = 12'b001110100111;
		12'b010000101010: color_data = 12'b001110100111;
		12'b010000110110: color_data = 12'b001110100111;
		12'b010000110111: color_data = 12'b001110100111;
		12'b010000111000: color_data = 12'b001110100111;
		12'b010000111001: color_data = 12'b001110100111;
		12'b010000111010: color_data = 12'b001110100111;
		12'b010001000011: color_data = 12'b001110100111;
		12'b010001000100: color_data = 12'b001110100111;
		12'b010001000101: color_data = 12'b001110100111;
		12'b010001001000: color_data = 12'b001110100111;
		12'b010001001001: color_data = 12'b001110100111;
		12'b010001001010: color_data = 12'b001110100111;
		12'b010001010011: color_data = 12'b001110100111;
		12'b010001010100: color_data = 12'b001110100111;
		12'b010001010101: color_data = 12'b001110100111;
		12'b010001011000: color_data = 12'b001110100111;
		12'b010001011001: color_data = 12'b001110100111;
		12'b010001011010: color_data = 12'b001110100111;
		12'b010001100000: color_data = 12'b001110100111;
		12'b010001100001: color_data = 12'b001110100111;
		12'b010001100010: color_data = 12'b001110100111;
		12'b010001101000: color_data = 12'b001110100111;
		12'b010001101001: color_data = 12'b001110100111;
		12'b010001101010: color_data = 12'b001110100111;
		12'b010001110000: color_data = 12'b001110100111;
		12'b010001110001: color_data = 12'b001110100111;
		12'b010001110010: color_data = 12'b001110100111;
		12'b010001111000: color_data = 12'b001110100111;
		12'b010001111001: color_data = 12'b001110100111;
		12'b010001111010: color_data = 12'b001110100111;
		12'b010010000000: color_data = 12'b001110100111;
		12'b010010000001: color_data = 12'b001110100111;
		12'b010010000010: color_data = 12'b001110100111;
		12'b010010000011: color_data = 12'b001110100111;
		12'b010010000100: color_data = 12'b001110100111;
		12'b010010000101: color_data = 12'b001110100111;
		12'b010010000110: color_data = 12'b001110100111;
		12'b010010000111: color_data = 12'b001110100111;
		12'b010010001000: color_data = 12'b001110100111;
		12'b010010001001: color_data = 12'b001110100111;
		12'b010010001010: color_data = 12'b001110100111;
		12'b010010001011: color_data = 12'b001110100111;
		12'b010010001100: color_data = 12'b001110100111;
		12'b010010010000: color_data = 12'b001110100111;
		12'b010010010001: color_data = 12'b001110100111;
		12'b010010010010: color_data = 12'b001110100111;
		12'b010010010011: color_data = 12'b001110100111;
		12'b010010010100: color_data = 12'b001110100111;
		12'b010010010101: color_data = 12'b001110100111;
		12'b010010010110: color_data = 12'b001110100111;
		12'b010010010111: color_data = 12'b001110100111;
		12'b010010011000: color_data = 12'b001110100111;
		12'b010010011001: color_data = 12'b001110100111;
		12'b010010011010: color_data = 12'b001110100111;
		12'b010010011011: color_data = 12'b001110100111;
		12'b010010011100: color_data = 12'b001110100111;
		12'b010010101000: color_data = 12'b001110100111;
		12'b010010101001: color_data = 12'b001110100111;
		12'b010010101010: color_data = 12'b001110100111;
		12'b010010111000: color_data = 12'b001110100111;
		12'b010010111001: color_data = 12'b001110100111;
		12'b010010111010: color_data = 12'b001110100111;
		12'b010011001000: color_data = 12'b001110100111;
		12'b010011001001: color_data = 12'b001110100111;
		12'b010011001010: color_data = 12'b001110100111;
		12'b010011011000: color_data = 12'b001110100111;
		12'b010011011001: color_data = 12'b001110100111;
		12'b010011011010: color_data = 12'b001110100111;
        12'b010100000000: color_data = 12'b001110100111;
		12'b010100000001: color_data = 12'b001110100111;
		12'b010100000010: color_data = 12'b001110100111;
		12'b010100000011: color_data = 12'b001110100111;
		12'b010100000100: color_data = 12'b001110100111;
		12'b010100000101: color_data = 12'b001110100111;
		12'b010100000110: color_data = 12'b001110100111;
		12'b010100000111: color_data = 12'b001110100111;
		12'b010100001000: color_data = 12'b001110100111;
		12'b010100001001: color_data = 12'b001110100111;
		12'b010100001010: color_data = 12'b001110100111;
		12'b010100001011: color_data = 12'b001110100111;
		12'b010100001100: color_data = 12'b001110100111;
		12'b010100010000: color_data = 12'b001110100111;
		12'b010100010001: color_data = 12'b001110100111;
		12'b010100010010: color_data = 12'b001110100111;
		12'b010100010011: color_data = 12'b001110100111;
		12'b010100010100: color_data = 12'b001110100111;
		12'b010100010101: color_data = 12'b001110100111;
		12'b010100010110: color_data = 12'b001110100111;
		12'b010100010111: color_data = 12'b001110100111;
		12'b010100011000: color_data = 12'b001110100111;
		12'b010100011001: color_data = 12'b001110100111;
		12'b010100011010: color_data = 12'b001110100111;
		12'b010100011011: color_data = 12'b001110100111;
		12'b010100011100: color_data = 12'b001110100111;
		12'b010100100000: color_data = 12'b001110100111;
		12'b010100100001: color_data = 12'b001110100111;
		12'b010100100010: color_data = 12'b001110100111;
		12'b010100110000: color_data = 12'b001110100111;
		12'b010100110001: color_data = 12'b001110100111;
		12'b010100110010: color_data = 12'b001110100111;
		12'b010101000000: color_data = 12'b001110100111;
		12'b010101000001: color_data = 12'b001110100111;
		12'b010101000010: color_data = 12'b001110100111;
		12'b010101000011: color_data = 12'b001110100111;
		12'b010101000100: color_data = 12'b001110100111;
		12'b010101000101: color_data = 12'b001110100111;
		12'b010101000110: color_data = 12'b001110100111;
		12'b010101000111: color_data = 12'b001110100111;
		12'b010101001000: color_data = 12'b001110100111;
		12'b010101001001: color_data = 12'b001110100111;
		12'b010101001010: color_data = 12'b001110100111;
		12'b010101010000: color_data = 12'b001110100111;
		12'b010101010001: color_data = 12'b001110100111;
		12'b010101010010: color_data = 12'b001110100111;
		12'b010101010011: color_data = 12'b001110100111;
		12'b010101010100: color_data = 12'b001110100111;
		12'b010101010101: color_data = 12'b001110100111;
		12'b010101010110: color_data = 12'b001110100111;
		12'b010101010111: color_data = 12'b001110100111;
		12'b010101011000: color_data = 12'b001110100111;
		12'b010101011001: color_data = 12'b001110100111;
		12'b010101011010: color_data = 12'b001110100111;
		12'b010101100110: color_data = 12'b001110100111;
		12'b010101100111: color_data = 12'b001110100111;
		12'b010101101011: color_data = 12'b001110100111;
		12'b010101101100: color_data = 12'b001110100111;
		12'b010101110110: color_data = 12'b001110100111;
		12'b010101110111: color_data = 12'b001110100111;
		12'b010101111011: color_data = 12'b001110100111;
		12'b010101111100: color_data = 12'b001110100111;
		12'b010110001011: color_data = 12'b001110100111;
		12'b010110001100: color_data = 12'b001110100111;
		12'b010110011011: color_data = 12'b001110100111;
		12'b010110011100: color_data = 12'b001110100111;
		12'b010110100110: color_data = 12'b001110100111;
		12'b010110100111: color_data = 12'b001110100111;
		12'b010110101011: color_data = 12'b001110100111;
		12'b010110101100: color_data = 12'b001110100111;
		12'b010110110110: color_data = 12'b001110100111;
		12'b010110110111: color_data = 12'b001110100111;
		12'b010110111011: color_data = 12'b001110100111;
		12'b010110111100: color_data = 12'b001110100111;
		12'b010111000000: color_data = 12'b001110100111;
		12'b010111000001: color_data = 12'b001110100111;
		12'b010111000010: color_data = 12'b001110100111;
		12'b010111000011: color_data = 12'b001110100111;
		12'b010111000100: color_data = 12'b001110100111;
		12'b010111000101: color_data = 12'b001110100111;
		12'b010111000110: color_data = 12'b001110100111;
		12'b010111000111: color_data = 12'b001110100111;
		12'b010111001000: color_data = 12'b001110100111;
		12'b010111001001: color_data = 12'b001110100111;
		12'b010111001010: color_data = 12'b001110100111;
		12'b010111010000: color_data = 12'b001110100111;
		12'b010111010001: color_data = 12'b001110100111;
		12'b010111010010: color_data = 12'b001110100111;
		12'b010111010011: color_data = 12'b001110100111;
		12'b010111010100: color_data = 12'b001110100111;
		12'b010111010101: color_data = 12'b001110100111;
		12'b010111010110: color_data = 12'b001110100111;
		12'b010111010111: color_data = 12'b001110100111;
		12'b010111011000: color_data = 12'b001110100111;
		12'b010111011001: color_data = 12'b001110100111;
		12'b010111011010: color_data = 12'b001110100111;
        12'b011000000011: color_data = 12'b001110100111;
		12'b011000000100: color_data = 12'b001110100111;
		12'b011000000101: color_data = 12'b001110100111;
		12'b011000000110: color_data = 12'b001110100111;
		12'b011000000111: color_data = 12'b001110100111;
		12'b011000001000: color_data = 12'b001110100111;
		12'b011000001001: color_data = 12'b001110100111;
		12'b011000001010: color_data = 12'b001110100111;
		12'b011000010011: color_data = 12'b001110100111;
		12'b011000010100: color_data = 12'b001110100111;
		12'b011000010101: color_data = 12'b001110100111;
		12'b011000010110: color_data = 12'b001110100111;
		12'b011000010111: color_data = 12'b001110100111;
		12'b011000011000: color_data = 12'b001110100111;
		12'b011000011001: color_data = 12'b001110100111;
		12'b011000011010: color_data = 12'b001110100111;
		12'b011000100000: color_data = 12'b001110100111;
		12'b011000100001: color_data = 12'b001110100111;
		12'b011000100010: color_data = 12'b001110100111;
		12'b011000110000: color_data = 12'b001110100111;
		12'b011000110001: color_data = 12'b001110100111;
		12'b011000110010: color_data = 12'b001110100111;
		12'b011001000000: color_data = 12'b001110100111;
		12'b011001000001: color_data = 12'b001110100111;
		12'b011001000010: color_data = 12'b001110100111;
		12'b011001000011: color_data = 12'b001110100111;
		12'b011001000100: color_data = 12'b001110100111;
		12'b011001000101: color_data = 12'b001110100111;
		12'b011001000110: color_data = 12'b001110100111;
		12'b011001000111: color_data = 12'b001110100111;
		12'b011001001000: color_data = 12'b001110100111;
		12'b011001001001: color_data = 12'b001110100111;
		12'b011001001010: color_data = 12'b001110100111;
		12'b011001010000: color_data = 12'b001110100111;
		12'b011001010001: color_data = 12'b001110100111;
		12'b011001010010: color_data = 12'b001110100111;
		12'b011001010011: color_data = 12'b001110100111;
		12'b011001010100: color_data = 12'b001110100111;
		12'b011001010101: color_data = 12'b001110100111;
		12'b011001010110: color_data = 12'b001110100111;
		12'b011001010111: color_data = 12'b001110100111;
		12'b011001011000: color_data = 12'b001110100111;
		12'b011001011001: color_data = 12'b001110100111;
		12'b011001011010: color_data = 12'b001110100111;
		12'b011001100000: color_data = 12'b001110100111;
		12'b011001100001: color_data = 12'b001110100111;
		12'b011001100010: color_data = 12'b001110100111;
		12'b011001101011: color_data = 12'b001110100111;
		12'b011001101100: color_data = 12'b001110100111;
		12'b011001110000: color_data = 12'b001110100111;
		12'b011001110001: color_data = 12'b001110100111;
		12'b011001110010: color_data = 12'b001110100111;
		12'b011001111011: color_data = 12'b001110100111;
		12'b011001111100: color_data = 12'b001110100111;
		12'b011010000000: color_data = 12'b001110100111;
		12'b011010000001: color_data = 12'b001110100111;
		12'b011010000010: color_data = 12'b001110100111;
		12'b011010001011: color_data = 12'b001110100111;
		12'b011010001100: color_data = 12'b001110100111;
		12'b011010010000: color_data = 12'b001110100111;
		12'b011010010001: color_data = 12'b001110100111;
		12'b011010010010: color_data = 12'b001110100111;
		12'b011010011011: color_data = 12'b001110100111;
		12'b011010011100: color_data = 12'b001110100111;
		12'b011010100000: color_data = 12'b001110100111;
		12'b011010100001: color_data = 12'b001110100111;
		12'b011010100010: color_data = 12'b001110100111;
		12'b011010101011: color_data = 12'b001110100111;
		12'b011010101100: color_data = 12'b001110100111;
		12'b011010110000: color_data = 12'b001110100111;
		12'b011010110001: color_data = 12'b001110100111;
		12'b011010110010: color_data = 12'b001110100111;
		12'b011010111011: color_data = 12'b001110100111;
		12'b011010111100: color_data = 12'b001110100111;
		12'b011011000011: color_data = 12'b001110100111;
		12'b011011000100: color_data = 12'b001110100111;
		12'b011011000101: color_data = 12'b001110100111;
		12'b011011000110: color_data = 12'b001110100111;
		12'b011011000111: color_data = 12'b001110100111;
		12'b011011001000: color_data = 12'b001110100111;
		12'b011011001001: color_data = 12'b001110100111;
		12'b011011001010: color_data = 12'b001110100111;
		12'b011011010011: color_data = 12'b001110100111;
		12'b011011010100: color_data = 12'b001110100111;
		12'b011011010101: color_data = 12'b001110100111;
		12'b011011010110: color_data = 12'b001110100111;
		12'b011011010111: color_data = 12'b001110100111;
		12'b011011011000: color_data = 12'b001110100111;
		12'b011011011001: color_data = 12'b001110100111;
		12'b011011011010: color_data = 12'b001110100111;
        12'b011100000000: color_data = 12'b001110100111;
		12'b011100000001: color_data = 12'b001110100111;
		12'b011100000010: color_data = 12'b001110100111;
		12'b011100000011: color_data = 12'b001110100111;
		12'b011100000100: color_data = 12'b001110100111;
		12'b011100000101: color_data = 12'b001110100111;
		12'b011100000110: color_data = 12'b001110100111;
		12'b011100000111: color_data = 12'b001110100111;
		12'b011100001000: color_data = 12'b001110100111;
		12'b011100001001: color_data = 12'b001110100111;
		12'b011100001010: color_data = 12'b001110100111;
		12'b011100001011: color_data = 12'b001110100111;
		12'b011100001100: color_data = 12'b001110100111;
		12'b011100010000: color_data = 12'b001110100111;
		12'b011100010001: color_data = 12'b001110100111;
		12'b011100010010: color_data = 12'b001110100111;
		12'b011100010011: color_data = 12'b001110100111;
		12'b011100010100: color_data = 12'b001110100111;
		12'b011100010101: color_data = 12'b001110100111;
		12'b011100010110: color_data = 12'b001110100111;
		12'b011100010111: color_data = 12'b001110100111;
		12'b011100011000: color_data = 12'b001110100111;
		12'b011100011001: color_data = 12'b001110100111;
		12'b011100011010: color_data = 12'b001110100111;
		12'b011100011011: color_data = 12'b001110100111;
		12'b011100011100: color_data = 12'b001110100111;
		12'b011100101011: color_data = 12'b001110100111;
		12'b011100101100: color_data = 12'b001110100111;
		12'b011100111011: color_data = 12'b001110100111;
		12'b011100111100: color_data = 12'b001110100111;
		12'b011101001011: color_data = 12'b001110100111;
		12'b011101001100: color_data = 12'b001110100111;
		12'b011101011011: color_data = 12'b001110100111;
		12'b011101011100: color_data = 12'b001110100111;
		12'b011101101000: color_data = 12'b001110100111;
		12'b011101101001: color_data = 12'b001110100111;
		12'b011101101010: color_data = 12'b001110100111;
		12'b011101111000: color_data = 12'b001110100111;
		12'b011101111001: color_data = 12'b001110100111;
		12'b011101111010: color_data = 12'b001110100111;
		12'b011110001000: color_data = 12'b001110100111;
		12'b011110001001: color_data = 12'b001110100111;
		12'b011110001010: color_data = 12'b001110100111;
		12'b011110011000: color_data = 12'b001110100111;
		12'b011110011001: color_data = 12'b001110100111;
		12'b011110011010: color_data = 12'b001110100111;
		12'b011110100110: color_data = 12'b001110100111;
		12'b011110100111: color_data = 12'b001110100111;
		12'b011110110110: color_data = 12'b001110100111;
		12'b011110110111: color_data = 12'b001110100111;
		12'b011111000110: color_data = 12'b001110100111;
		12'b011111000111: color_data = 12'b001110100111;
		12'b011111010110: color_data = 12'b001110100111;
		12'b011111010111: color_data = 12'b001110100111;
        12'b100000000011: color_data = 12'b001110100111;
		12'b100000000100: color_data = 12'b001110100111;
		12'b100000000101: color_data = 12'b001110100111;
		12'b100000000110: color_data = 12'b001110100111;
		12'b100000000111: color_data = 12'b001110100111;
		12'b100000001000: color_data = 12'b001110100111;
		12'b100000001001: color_data = 12'b001110100111;
		12'b100000001010: color_data = 12'b001110100111;
		12'b100000010011: color_data = 12'b001110100111;
		12'b100000010100: color_data = 12'b001110100111;
		12'b100000010101: color_data = 12'b001110100111;
		12'b100000010110: color_data = 12'b001110100111;
		12'b100000010111: color_data = 12'b001110100111;
		12'b100000011000: color_data = 12'b001110100111;
		12'b100000011001: color_data = 12'b001110100111;
		12'b100000011010: color_data = 12'b001110100111;
		12'b100000100000: color_data = 12'b001110100111;
		12'b100000100001: color_data = 12'b001110100111;
		12'b100000100010: color_data = 12'b001110100111;
		12'b100000101011: color_data = 12'b001110100111;
		12'b100000101100: color_data = 12'b001110100111;
		12'b100000110000: color_data = 12'b001110100111;
		12'b100000110001: color_data = 12'b001110100111;
		12'b100000110010: color_data = 12'b001110100111;
		12'b100000111011: color_data = 12'b001110100111;
		12'b100000111100: color_data = 12'b001110100111;
		12'b100001000000: color_data = 12'b001110100111;
		12'b100001000001: color_data = 12'b001110100111;
		12'b100001000010: color_data = 12'b001110100111;
		12'b100001001011: color_data = 12'b001110100111;
		12'b100001001100: color_data = 12'b001110100111;
		12'b100001010000: color_data = 12'b001110100111;
		12'b100001010001: color_data = 12'b001110100111;
		12'b100001010010: color_data = 12'b001110100111;
		12'b100001011011: color_data = 12'b001110100111;
		12'b100001011100: color_data = 12'b001110100111;
		12'b100001100011: color_data = 12'b001110100111;
		12'b100001100100: color_data = 12'b001110100111;
		12'b100001100101: color_data = 12'b001110100111;
		12'b100001100110: color_data = 12'b001110100111;
		12'b100001100111: color_data = 12'b001110100111;
		12'b100001101000: color_data = 12'b001110100111;
		12'b100001101001: color_data = 12'b001110100111;
		12'b100001101010: color_data = 12'b001110100111;
		12'b100001110011: color_data = 12'b001110100111;
		12'b100001110100: color_data = 12'b001110100111;
		12'b100001110101: color_data = 12'b001110100111;
		12'b100001110110: color_data = 12'b001110100111;
		12'b100001110111: color_data = 12'b001110100111;
		12'b100001111000: color_data = 12'b001110100111;
		12'b100001111001: color_data = 12'b001110100111;
		12'b100001111010: color_data = 12'b001110100111;
		12'b100010000000: color_data = 12'b001110100111;
		12'b100010000001: color_data = 12'b001110100111;
		12'b100010000010: color_data = 12'b001110100111;
		12'b100010001011: color_data = 12'b001110100111;
		12'b100010001100: color_data = 12'b001110100111;
		12'b100010010000: color_data = 12'b001110100111;
		12'b100010010001: color_data = 12'b001110100111;
		12'b100010010010: color_data = 12'b001110100111;
		12'b100010011011: color_data = 12'b001110100111;
		12'b100010011100: color_data = 12'b001110100111;
		12'b100010100000: color_data = 12'b001110100111;
		12'b100010100001: color_data = 12'b001110100111;
		12'b100010100010: color_data = 12'b001110100111;
		12'b100010101011: color_data = 12'b001110100111;
		12'b100010101100: color_data = 12'b001110100111;
		12'b100010110000: color_data = 12'b001110100111;
		12'b100010110001: color_data = 12'b001110100111;
		12'b100010110010: color_data = 12'b001110100111;
		12'b100010111011: color_data = 12'b001110100111;
		12'b100010111100: color_data = 12'b001110100111;
		12'b100011000011: color_data = 12'b001110100111;
		12'b100011000100: color_data = 12'b001110100111;
		12'b100011000101: color_data = 12'b001110100111;
		12'b100011000110: color_data = 12'b001110100111;
		12'b100011000111: color_data = 12'b001110100111;
		12'b100011001000: color_data = 12'b001110100111;
		12'b100011001001: color_data = 12'b001110100111;
		12'b100011001010: color_data = 12'b001110100111;
		12'b100011010011: color_data = 12'b001110100111;
		12'b100011010100: color_data = 12'b001110100111;
		12'b100011010101: color_data = 12'b001110100111;
		12'b100011010110: color_data = 12'b001110100111;
		12'b100011010111: color_data = 12'b001110100111;
		12'b100011011000: color_data = 12'b001110100111;
		12'b100011011001: color_data = 12'b001110100111;
		12'b100011011010: color_data = 12'b001110100111;
        12'b100100000011: color_data = 12'b001110100111;
		12'b100100000100: color_data = 12'b001110100111;
		12'b100100000101: color_data = 12'b001110100111;
		12'b100100000110: color_data = 12'b001110100111;
		12'b100100000111: color_data = 12'b001110100111;
		12'b100100001000: color_data = 12'b001110100111;
		12'b100100001001: color_data = 12'b001110100111;
		12'b100100001010: color_data = 12'b001110100111;
		12'b100100010011: color_data = 12'b001110100111;
		12'b100100010100: color_data = 12'b001110100111;
		12'b100100010101: color_data = 12'b001110100111;
		12'b100100010110: color_data = 12'b001110100111;
		12'b100100010111: color_data = 12'b001110100111;
		12'b100100011000: color_data = 12'b001110100111;
		12'b100100011001: color_data = 12'b001110100111;
		12'b100100011010: color_data = 12'b001110100111;
		12'b100100100000: color_data = 12'b001110100111;
		12'b100100100001: color_data = 12'b001110100111;
		12'b100100100010: color_data = 12'b001110100111;
		12'b100100101011: color_data = 12'b001110100111;
		12'b100100101100: color_data = 12'b001110100111;
		12'b100100110000: color_data = 12'b001110100111;
		12'b100100110001: color_data = 12'b001110100111;
		12'b100100110010: color_data = 12'b001110100111;
		12'b100100111011: color_data = 12'b001110100111;
		12'b100100111100: color_data = 12'b001110100111;
		12'b100101000000: color_data = 12'b001110100111;
		12'b100101000001: color_data = 12'b001110100111;
		12'b100101000010: color_data = 12'b001110100111;
		12'b100101001011: color_data = 12'b001110100111;
		12'b100101001100: color_data = 12'b001110100111;
		12'b100101010000: color_data = 12'b001110100111;
		12'b100101010001: color_data = 12'b001110100111;
		12'b100101010010: color_data = 12'b001110100111;
		12'b100101011011: color_data = 12'b001110100111;
		12'b100101011100: color_data = 12'b001110100111;
		12'b100101100000: color_data = 12'b001110100111;
		12'b100101100001: color_data = 12'b001110100111;
		12'b100101100010: color_data = 12'b001110100111;
		12'b100101101011: color_data = 12'b001110100111;
		12'b100101101100: color_data = 12'b001110100111;
		12'b100101110000: color_data = 12'b001110100111;
		12'b100101110001: color_data = 12'b001110100111;
		12'b100101110010: color_data = 12'b001110100111;
		12'b100101111011: color_data = 12'b001110100111;
		12'b100101111100: color_data = 12'b001110100111;
		12'b100110000011: color_data = 12'b001110100111;
		12'b100110000100: color_data = 12'b001110100111;
		12'b100110000101: color_data = 12'b001110100111;
		12'b100110000110: color_data = 12'b001110100111;
		12'b100110000111: color_data = 12'b001110100111;
		12'b100110001000: color_data = 12'b001110100111;
		12'b100110001001: color_data = 12'b001110100111;
		12'b100110001010: color_data = 12'b001110100111;
		12'b100110001011: color_data = 12'b001110100111;
		12'b100110001100: color_data = 12'b001110100111;
		12'b100110010011: color_data = 12'b001110100111;
		12'b100110010100: color_data = 12'b001110100111;
		12'b100110010101: color_data = 12'b001110100111;
		12'b100110010110: color_data = 12'b001110100111;
		12'b100110010111: color_data = 12'b001110100111;
		12'b100110011000: color_data = 12'b001110100111;
		12'b100110011001: color_data = 12'b001110100111;
		12'b100110011010: color_data = 12'b001110100111;
		12'b100110011011: color_data = 12'b001110100111;
		12'b100110011100: color_data = 12'b001110100111;
		12'b100110101011: color_data = 12'b001110100111;
		12'b100110101100: color_data = 12'b001110100111;
		12'b100110111011: color_data = 12'b001110100111;
		12'b100110111100: color_data = 12'b001110100111;
		12'b100111000011: color_data = 12'b001110100111;
		12'b100111000100: color_data = 12'b001110100111;
		12'b100111000101: color_data = 12'b001110100111;
		12'b100111000110: color_data = 12'b001110100111;
		12'b100111000111: color_data = 12'b001110100111;
		12'b100111001000: color_data = 12'b001110100111;
		12'b100111001001: color_data = 12'b001110100111;
		12'b100111001010: color_data = 12'b001110100111;
		12'b100111010011: color_data = 12'b001110100111;
		12'b100111010100: color_data = 12'b001110100111;
		12'b100111010101: color_data = 12'b001110100111;
		12'b100111010110: color_data = 12'b001110100111;
		12'b100111010111: color_data = 12'b001110100111;
		12'b100111011000: color_data = 12'b001110100111;
		12'b100111011001: color_data = 12'b001110100111;
		12'b100111011010: color_data = 12'b001110100111;
		default: color_data = 12'b000000000000;
	endcase
endmodule
