`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.01.2025 14:29:31
// Design Name: 
// Module Name: continue_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module continue_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		13'b0000000110010: color_data = 12'b001110100111;
		13'b0000000110011: color_data = 12'b001110100111;
		13'b0000001000000: color_data = 12'b001110100111;
		13'b0000001000001: color_data = 12'b001110100111;
		13'b0000001011010: color_data = 12'b001110100111;
		13'b0000001011011: color_data = 12'b001110100111;
		13'b0000001011100: color_data = 12'b001110100111;
		13'b0000001100100: color_data = 12'b001110100111;
		13'b0000001100101: color_data = 12'b001110100111;
		13'b0000001100110: color_data = 12'b001110100111;
		13'b0000001100111: color_data = 12'b001110100111;
		13'b0000001101000: color_data = 12'b001110100111;
		13'b0000100000011: color_data = 12'b001110100111;
		13'b0000100000100: color_data = 12'b001110100111;
		13'b0000100000101: color_data = 12'b001110100111;
		13'b0000100000110: color_data = 12'b001110100111;
		13'b0000100000111: color_data = 12'b001110100111;
		13'b0000100001000: color_data = 12'b001110100111;
		13'b0000100001001: color_data = 12'b001110100111;
		13'b0000100001010: color_data = 12'b001110100111;
		13'b0000100001011: color_data = 12'b001110100111;
		13'b0000100010011: color_data = 12'b001110100111;
		13'b0000100010100: color_data = 12'b001110100111;
		13'b0000100010101: color_data = 12'b001110100111;
		13'b0000100010110: color_data = 12'b001110100111;
		13'b0000100010111: color_data = 12'b001110100111;
		13'b0000100011000: color_data = 12'b001110100111;
		13'b0000100011001: color_data = 12'b001110100111;
		13'b0000100011010: color_data = 12'b001110100111;
		13'b0000100011011: color_data = 12'b001110100111;
		13'b0000100100000: color_data = 12'b001110100111;
		13'b0000100100001: color_data = 12'b001110100111;
		13'b0000100100010: color_data = 12'b001110100111;
		13'b0000100100011: color_data = 12'b001110100111;
		13'b0000100101101: color_data = 12'b001110100111;
		13'b0000100101110: color_data = 12'b001110100111;
		13'b0000100101111: color_data = 12'b001110100111;
		13'b0000100110000: color_data = 12'b001110100111;
		13'b0000100110010: color_data = 12'b001110100111;
		13'b0000100110011: color_data = 12'b001110100111;
		13'b0000100110100: color_data = 12'b001110100111;
		13'b0000100110101: color_data = 12'b001110100111;
		13'b0000100110110: color_data = 12'b001110100111;
		13'b0000100110111: color_data = 12'b001110100111;
		13'b0000100111000: color_data = 12'b001110100111;
		13'b0000100111001: color_data = 12'b001110100111;
		13'b0000100111010: color_data = 12'b001110100111;
		13'b0000100111011: color_data = 12'b001110100111;
		13'b0000100111100: color_data = 12'b001110100111;
		13'b0000100111101: color_data = 12'b001110100111;
		13'b0000100111110: color_data = 12'b001110100111;
		13'b0000100111111: color_data = 12'b001110100111;
		13'b0000101000000: color_data = 12'b001110100111;
		13'b0000101000001: color_data = 12'b001110100111;
		13'b0000101000011: color_data = 12'b001110100111;
		13'b0000101000100: color_data = 12'b001110100111;
		13'b0000101000101: color_data = 12'b001110100111;
		13'b0000101000110: color_data = 12'b001110100111;
		13'b0000101001000: color_data = 12'b001110100111;
		13'b0000101001001: color_data = 12'b001110100111;
		13'b0000101001010: color_data = 12'b001110100111;
		13'b0000101001011: color_data = 12'b001110100111;
		13'b0000101010101: color_data = 12'b001110100111;
		13'b0000101010110: color_data = 12'b001110100111;
		13'b0000101010111: color_data = 12'b001110100111;
		13'b0000101011000: color_data = 12'b001110100111;
		13'b0000101011010: color_data = 12'b001110100111;
		13'b0000101011011: color_data = 12'b001110100111;
		13'b0000101011100: color_data = 12'b001110100111;
		13'b0000101100100: color_data = 12'b001110100111;
		13'b0000101100101: color_data = 12'b001110100111;
		13'b0000101100110: color_data = 12'b001110100111;
		13'b0000101101000: color_data = 12'b001110100111;
		13'b0000101101010: color_data = 12'b001110100111;
		13'b0000101101011: color_data = 12'b001110100111;
		13'b0000101101100: color_data = 12'b001110100111;
		13'b0000101101101: color_data = 12'b001110100111;
		13'b0000101101110: color_data = 12'b001110100111;
		13'b0000101101111: color_data = 12'b001110100111;
		13'b0000101110000: color_data = 12'b001110100111;
		13'b0000101110001: color_data = 12'b001110100111;
		13'b0000101110010: color_data = 12'b001110100111;
		13'b0000101110011: color_data = 12'b001110100111;
		13'b0000101110100: color_data = 12'b001110100111;
		13'b0000101110101: color_data = 12'b001110100111;
		13'b0000101110110: color_data = 12'b001110100111;
		13'b0000101111100: color_data = 12'b001110100111;
		13'b0000101111101: color_data = 12'b001110100111;
		13'b0000101111110: color_data = 12'b001110100111;
		13'b0000101111111: color_data = 12'b001110100111;
		13'b0000110000000: color_data = 12'b001110100111;
		13'b0000110000001: color_data = 12'b001110100111;
		13'b0000110000010: color_data = 12'b001110100111;
		13'b0000110000011: color_data = 12'b001110100111;
		13'b0000110000100: color_data = 12'b001110100111;
		13'b0001000000010: color_data = 12'b001110100111;
		13'b0001000000011: color_data = 12'b001110100111;
		13'b0001000000100: color_data = 12'b001110100111;
		13'b0001000000101: color_data = 12'b001110100111;
		13'b0001000000110: color_data = 12'b001110100111;
		13'b0001000000111: color_data = 12'b001110100111;
		13'b0001000001000: color_data = 12'b001110100111;
		13'b0001000001001: color_data = 12'b001110100111;
		13'b0001000001010: color_data = 12'b001110100111;
		13'b0001000001011: color_data = 12'b001110100111;
		13'b0001000001100: color_data = 12'b001110100111;
		13'b0001000010010: color_data = 12'b001110100111;
		13'b0001000010011: color_data = 12'b001110100111;
		13'b0001000010100: color_data = 12'b001110100111;
		13'b0001000010101: color_data = 12'b001110100111;
		13'b0001000010110: color_data = 12'b001110100111;
		13'b0001000010111: color_data = 12'b001110100111;
		13'b0001000011000: color_data = 12'b001110100111;
		13'b0001000011001: color_data = 12'b001110100111;
		13'b0001000011010: color_data = 12'b001110100111;
		13'b0001000011011: color_data = 12'b001110100111;
		13'b0001000011100: color_data = 12'b001110100111;
		13'b0001000100000: color_data = 12'b001110100111;
		13'b0001000100001: color_data = 12'b001110100111;
		13'b0001000100010: color_data = 12'b001110100111;
		13'b0001000100011: color_data = 12'b001110100111;
		13'b0001000101101: color_data = 12'b001110100111;
		13'b0001000101110: color_data = 12'b001110100111;
		13'b0001000101111: color_data = 12'b001110100111;
		13'b0001000110000: color_data = 12'b001110100111;
		13'b0001000110010: color_data = 12'b001110100111;
		13'b0001000110011: color_data = 12'b001110100111;
		13'b0001000110100: color_data = 12'b001110100111;
		13'b0001000110101: color_data = 12'b001110100111;
		13'b0001000110110: color_data = 12'b001110100111;
		13'b0001000110111: color_data = 12'b001110100111;
		13'b0001000111000: color_data = 12'b001110100111;
		13'b0001000111001: color_data = 12'b001110100111;
		13'b0001000111010: color_data = 12'b001110100111;
		13'b0001000111011: color_data = 12'b001110100111;
		13'b0001000111100: color_data = 12'b001110100111;
		13'b0001000111101: color_data = 12'b001110100111;
		13'b0001000111110: color_data = 12'b001110100111;
		13'b0001000111111: color_data = 12'b001110100111;
		13'b0001001000000: color_data = 12'b001110100111;
		13'b0001001000001: color_data = 12'b001110100111;
		13'b0001001000011: color_data = 12'b001110100111;
		13'b0001001000100: color_data = 12'b001110100111;
		13'b0001001000101: color_data = 12'b001110100111;
		13'b0001001000110: color_data = 12'b001110100111;
		13'b0001001001000: color_data = 12'b001110100111;
		13'b0001001001001: color_data = 12'b001110100111;
		13'b0001001001010: color_data = 12'b001110100111;
		13'b0001001001011: color_data = 12'b001110100111;
		13'b0001001010101: color_data = 12'b001110100111;
		13'b0001001010110: color_data = 12'b001110100111;
		13'b0001001010111: color_data = 12'b001110100111;
		13'b0001001011000: color_data = 12'b001110100111;
		13'b0001001011010: color_data = 12'b001110100111;
		13'b0001001011011: color_data = 12'b001110100111;
		13'b0001001011100: color_data = 12'b001110100111;
		13'b0001001100100: color_data = 12'b001110100111;
		13'b0001001100101: color_data = 12'b001110100111;
		13'b0001001100110: color_data = 12'b001110100111;
		13'b0001001101000: color_data = 12'b001110100111;
		13'b0001001101010: color_data = 12'b001110100111;
		13'b0001001101011: color_data = 12'b001110100111;
		13'b0001001101100: color_data = 12'b001110100111;
		13'b0001001101101: color_data = 12'b001110100111;
		13'b0001001101110: color_data = 12'b001110100111;
		13'b0001001101111: color_data = 12'b001110100111;
		13'b0001001110000: color_data = 12'b001110100111;
		13'b0001001110001: color_data = 12'b001110100111;
		13'b0001001110010: color_data = 12'b001110100111;
		13'b0001001110011: color_data = 12'b001110100111;
		13'b0001001110100: color_data = 12'b001110100111;
		13'b0001001110101: color_data = 12'b001110100111;
		13'b0001001110110: color_data = 12'b001110100111;
		13'b0001001111011: color_data = 12'b001110100111;
		13'b0001001111100: color_data = 12'b001110100111;
		13'b0001001111101: color_data = 12'b001110100111;
		13'b0001001111110: color_data = 12'b001110100111;
		13'b0001001111111: color_data = 12'b001110100111;
		13'b0001010000000: color_data = 12'b001110100111;
		13'b0001010000001: color_data = 12'b001110100111;
		13'b0001010000010: color_data = 12'b001110100111;
		13'b0001010000011: color_data = 12'b001110100111;
		13'b0001010000100: color_data = 12'b001110100111;
		13'b0001010000101: color_data = 12'b001110100111;
		13'b0001100000001: color_data = 12'b001110100111;
		13'b0001100000010: color_data = 12'b001110100111;
		13'b0001100000011: color_data = 12'b001110100111;
		13'b0001100000100: color_data = 12'b001110100111;
		13'b0001100001010: color_data = 12'b001110100111;
		13'b0001100001011: color_data = 12'b001110100111;
		13'b0001100001100: color_data = 12'b001110100111;
		13'b0001100001101: color_data = 12'b001110100111;
		13'b0001100010001: color_data = 12'b001110100111;
		13'b0001100010010: color_data = 12'b001110100111;
		13'b0001100010011: color_data = 12'b001110100111;
		13'b0001100011010: color_data = 12'b001110100111;
		13'b0001100011011: color_data = 12'b001110100111;
		13'b0001100011100: color_data = 12'b001110100111;
		13'b0001100011101: color_data = 12'b001110100111;
		13'b0001100100000: color_data = 12'b001110100111;
		13'b0001100100001: color_data = 12'b001110100111;
		13'b0001100100010: color_data = 12'b001110100111;
		13'b0001100100011: color_data = 12'b001110100111;
		13'b0001100101101: color_data = 12'b001110100111;
		13'b0001100101110: color_data = 12'b001110100111;
		13'b0001100110000: color_data = 12'b001110100111;
		13'b0001100110010: color_data = 12'b001110100111;
		13'b0001100110011: color_data = 12'b001110100111;
		13'b0001100110100: color_data = 12'b001110100111;
		13'b0001100110101: color_data = 12'b001110100111;
		13'b0001100110110: color_data = 12'b001110100111;
		13'b0001100110111: color_data = 12'b001110100111;
		13'b0001100111000: color_data = 12'b001110100111;
		13'b0001100111001: color_data = 12'b001110100111;
		13'b0001100111010: color_data = 12'b001110100111;
		13'b0001100111011: color_data = 12'b001110100111;
		13'b0001100111100: color_data = 12'b001110100111;
		13'b0001100111101: color_data = 12'b001110100111;
		13'b0001100111110: color_data = 12'b001110100111;
		13'b0001100111111: color_data = 12'b001110100111;
		13'b0001101000000: color_data = 12'b001110100111;
		13'b0001101000001: color_data = 12'b001110100111;
		13'b0001101000011: color_data = 12'b001110100111;
		13'b0001101000100: color_data = 12'b001110100111;
		13'b0001101000110: color_data = 12'b001110100111;
		13'b0001101001000: color_data = 12'b001110100111;
		13'b0001101001001: color_data = 12'b001110100111;
		13'b0001101001010: color_data = 12'b001110100111;
		13'b0001101001011: color_data = 12'b001110100111;
		13'b0001101010101: color_data = 12'b001110100111;
		13'b0001101010110: color_data = 12'b001110100111;
		13'b0001101011000: color_data = 12'b001110100111;
		13'b0001101011010: color_data = 12'b001110100111;
		13'b0001101011011: color_data = 12'b001110100111;
		13'b0001101011100: color_data = 12'b001110100111;
		13'b0001101100100: color_data = 12'b001110100111;
		13'b0001101100101: color_data = 12'b001110100111;
		13'b0001101100110: color_data = 12'b001110100111;
		13'b0001101101000: color_data = 12'b001110100111;
		13'b0001101101010: color_data = 12'b001110100111;
		13'b0001101101011: color_data = 12'b001110100111;
		13'b0001101101101: color_data = 12'b001110100111;
		13'b0001101110100: color_data = 12'b001110100111;
		13'b0001101110101: color_data = 12'b001110100111;
		13'b0001101110110: color_data = 12'b001110100111;
		13'b0001101110111: color_data = 12'b001110100111;
		13'b0001101111010: color_data = 12'b001110100111;
		13'b0001101111011: color_data = 12'b001110100111;
		13'b0001101111100: color_data = 12'b001110100111;
		13'b0001110000011: color_data = 12'b001110100111;
		13'b0001110000100: color_data = 12'b001110100111;
		13'b0001110000101: color_data = 12'b001110100111;
		13'b0001110000110: color_data = 12'b001110100111;
		13'b0010000000001: color_data = 12'b001110100111;
		13'b0010000000010: color_data = 12'b001110100111;
		13'b0010000000011: color_data = 12'b001110100111;
		13'b0010000000100: color_data = 12'b001110100111;
		13'b0010000001011: color_data = 12'b001110100111;
		13'b0010000001100: color_data = 12'b001110100111;
		13'b0010000001101: color_data = 12'b001110100111;
		13'b0010000010000: color_data = 12'b001110100111;
		13'b0010000010001: color_data = 12'b001110100111;
		13'b0010000010010: color_data = 12'b001110100111;
		13'b0010000011010: color_data = 12'b001110100111;
		13'b0010000011100: color_data = 12'b001110100111;
		13'b0010000011101: color_data = 12'b001110100111;
		13'b0010000011110: color_data = 12'b001110100111;
		13'b0010000100000: color_data = 12'b001110100111;
		13'b0010000100001: color_data = 12'b001110100111;
		13'b0010000100010: color_data = 12'b001110100111;
		13'b0010000100011: color_data = 12'b001110100111;
		13'b0010000100100: color_data = 12'b001110100111;
		13'b0010000101101: color_data = 12'b001110100111;
		13'b0010000101110: color_data = 12'b001110100111;
		13'b0010000110000: color_data = 12'b001110100111;
		13'b0010000110010: color_data = 12'b001110100111;
		13'b0010000110011: color_data = 12'b001110100111;
		13'b0010000111000: color_data = 12'b001110100111;
		13'b0010000111001: color_data = 12'b001110100111;
		13'b0010000111010: color_data = 12'b001110100111;
		13'b0010000111100: color_data = 12'b001110100111;
		13'b0010001000000: color_data = 12'b001110100111;
		13'b0010001000001: color_data = 12'b001110100111;
		13'b0010001000011: color_data = 12'b001110100111;
		13'b0010001000100: color_data = 12'b001110100111;
		13'b0010001000110: color_data = 12'b001110100111;
		13'b0010001001000: color_data = 12'b001110100111;
		13'b0010001001001: color_data = 12'b001110100111;
		13'b0010001001010: color_data = 12'b001110100111;
		13'b0010001001011: color_data = 12'b001110100111;
		13'b0010001001100: color_data = 12'b001110100111;
		13'b0010001010101: color_data = 12'b001110100111;
		13'b0010001010110: color_data = 12'b001110100111;
		13'b0010001011000: color_data = 12'b001110100111;
		13'b0010001011010: color_data = 12'b001110100111;
		13'b0010001011011: color_data = 12'b001110100111;
		13'b0010001011100: color_data = 12'b001110100111;
		13'b0010001100100: color_data = 12'b001110100111;
		13'b0010001100101: color_data = 12'b001110100111;
		13'b0010001100110: color_data = 12'b001110100111;
		13'b0010001101000: color_data = 12'b001110100111;
		13'b0010001101010: color_data = 12'b001110100111;
		13'b0010001101011: color_data = 12'b001110100111;
		13'b0010001101101: color_data = 12'b001110100111;
		13'b0010001110101: color_data = 12'b001110100111;
		13'b0010001110110: color_data = 12'b001110100111;
		13'b0010001110111: color_data = 12'b001110100111;
		13'b0010001111001: color_data = 12'b001110100111;
		13'b0010001111010: color_data = 12'b001110100111;
		13'b0010001111011: color_data = 12'b001110100111;
		13'b0010010000011: color_data = 12'b001110100111;
		13'b0010010000101: color_data = 12'b001110100111;
		13'b0010010000110: color_data = 12'b001110100111;
		13'b0010010000111: color_data = 12'b001110100111;
		13'b0010100000000: color_data = 12'b001110100111;
		13'b0010100000001: color_data = 12'b001110100111;
		13'b0010100000010: color_data = 12'b001110100111;
		13'b0010100000100: color_data = 12'b001110100111;
		13'b0010100001100: color_data = 12'b001110100111;
		13'b0010100001101: color_data = 12'b001110100111;
		13'b0010100001110: color_data = 12'b001110100111;
		13'b0010100010000: color_data = 12'b001110100111;
		13'b0010100010001: color_data = 12'b001110100111;
		13'b0010100010010: color_data = 12'b001110100111;
		13'b0010100011010: color_data = 12'b001110100111;
		13'b0010100011100: color_data = 12'b001110100111;
		13'b0010100011101: color_data = 12'b001110100111;
		13'b0010100011110: color_data = 12'b001110100111;
		13'b0010100100000: color_data = 12'b001110100111;
		13'b0010100100001: color_data = 12'b001110100111;
		13'b0010100100010: color_data = 12'b001110100111;
		13'b0010100100011: color_data = 12'b001110100111;
		13'b0010100100100: color_data = 12'b001110100111;
		13'b0010100101101: color_data = 12'b001110100111;
		13'b0010100101110: color_data = 12'b001110100111;
		13'b0010100110000: color_data = 12'b001110100111;
		13'b0010100111000: color_data = 12'b001110100111;
		13'b0010100111001: color_data = 12'b001110100111;
		13'b0010100111010: color_data = 12'b001110100111;
		13'b0010100111100: color_data = 12'b001110100111;
		13'b0010101000011: color_data = 12'b001110100111;
		13'b0010101000100: color_data = 12'b001110100111;
		13'b0010101000110: color_data = 12'b001110100111;
		13'b0010101001000: color_data = 12'b001110100111;
		13'b0010101001001: color_data = 12'b001110100111;
		13'b0010101001010: color_data = 12'b001110100111;
		13'b0010101001011: color_data = 12'b001110100111;
		13'b0010101001100: color_data = 12'b001110100111;
		13'b0010101010101: color_data = 12'b001110100111;
		13'b0010101010110: color_data = 12'b001110100111;
		13'b0010101011000: color_data = 12'b001110100111;
		13'b0010101011010: color_data = 12'b001110100111;
		13'b0010101011011: color_data = 12'b001110100111;
		13'b0010101011100: color_data = 12'b001110100111;
		13'b0010101100100: color_data = 12'b001110100111;
		13'b0010101100101: color_data = 12'b001110100111;
		13'b0010101100110: color_data = 12'b001110100111;
		13'b0010101101000: color_data = 12'b001110100111;
		13'b0010101101010: color_data = 12'b001110100111;
		13'b0010101101011: color_data = 12'b001110100111;
		13'b0010101101101: color_data = 12'b001110100111;
		13'b0010101111001: color_data = 12'b001110100111;
		13'b0010101111010: color_data = 12'b001110100111;
		13'b0010101111011: color_data = 12'b001110100111;
		13'b0010110000011: color_data = 12'b001110100111;
		13'b0010110000101: color_data = 12'b001110100111;
		13'b0010110000110: color_data = 12'b001110100111;
		13'b0010110000111: color_data = 12'b001110100111;
		13'b0011000000000: color_data = 12'b001110100111;
		13'b0011000000001: color_data = 12'b001110100111;
		13'b0011000000010: color_data = 12'b001110100111;
		13'b0011000000100: color_data = 12'b001110100111;
		13'b0011000001100: color_data = 12'b001110100111;
		13'b0011000001101: color_data = 12'b001110100111;
		13'b0011000001110: color_data = 12'b001110100111;
		13'b0011000010000: color_data = 12'b001110100111;
		13'b0011000010001: color_data = 12'b001110100111;
		13'b0011000010010: color_data = 12'b001110100111;
		13'b0011000011010: color_data = 12'b001110100111;
		13'b0011000011100: color_data = 12'b001110100111;
		13'b0011000011101: color_data = 12'b001110100111;
		13'b0011000011110: color_data = 12'b001110100111;
		13'b0011000100000: color_data = 12'b001110100111;
		13'b0011000100001: color_data = 12'b001110100111;
		13'b0011000100011: color_data = 12'b001110100111;
		13'b0011000100100: color_data = 12'b001110100111;
		13'b0011000100101: color_data = 12'b001110100111;
		13'b0011000101101: color_data = 12'b001110100111;
		13'b0011000101110: color_data = 12'b001110100111;
		13'b0011000110000: color_data = 12'b001110100111;
		13'b0011000111000: color_data = 12'b001110100111;
		13'b0011000111001: color_data = 12'b001110100111;
		13'b0011000111010: color_data = 12'b001110100111;
		13'b0011000111100: color_data = 12'b001110100111;
		13'b0011001000011: color_data = 12'b001110100111;
		13'b0011001000100: color_data = 12'b001110100111;
		13'b0011001000110: color_data = 12'b001110100111;
		13'b0011001001000: color_data = 12'b001110100111;
		13'b0011001001001: color_data = 12'b001110100111;
		13'b0011001001011: color_data = 12'b001110100111;
		13'b0011001001100: color_data = 12'b001110100111;
		13'b0011001001101: color_data = 12'b001110100111;
		13'b0011001010101: color_data = 12'b001110100111;
		13'b0011001010110: color_data = 12'b001110100111;
		13'b0011001011000: color_data = 12'b001110100111;
		13'b0011001011010: color_data = 12'b001110100111;
		13'b0011001011011: color_data = 12'b001110100111;
		13'b0011001011100: color_data = 12'b001110100111;
		13'b0011001100100: color_data = 12'b001110100111;
		13'b0011001100101: color_data = 12'b001110100111;
		13'b0011001100110: color_data = 12'b001110100111;
		13'b0011001101000: color_data = 12'b001110100111;
		13'b0011001101010: color_data = 12'b001110100111;
		13'b0011001101011: color_data = 12'b001110100111;
		13'b0011001101101: color_data = 12'b001110100111;
		13'b0011001111001: color_data = 12'b001110100111;
		13'b0011001111010: color_data = 12'b001110100111;
		13'b0011001111011: color_data = 12'b001110100111;
		13'b0011010000011: color_data = 12'b001110100111;
		13'b0011010000101: color_data = 12'b001110100111;
		13'b0011010000110: color_data = 12'b001110100111;
		13'b0011010000111: color_data = 12'b001110100111;
		13'b0011100000000: color_data = 12'b001110100111;
		13'b0011100000001: color_data = 12'b001110100111;
		13'b0011100000010: color_data = 12'b001110100111;
		13'b0011100000100: color_data = 12'b001110100111;
		13'b0011100010000: color_data = 12'b001110100111;
		13'b0011100010001: color_data = 12'b001110100111;
		13'b0011100010010: color_data = 12'b001110100111;
		13'b0011100011010: color_data = 12'b001110100111;
		13'b0011100011100: color_data = 12'b001110100111;
		13'b0011100011101: color_data = 12'b001110100111;
		13'b0011100011110: color_data = 12'b001110100111;
		13'b0011100100000: color_data = 12'b001110100111;
		13'b0011100100001: color_data = 12'b001110100111;
		13'b0011100100011: color_data = 12'b001110100111;
		13'b0011100100100: color_data = 12'b001110100111;
		13'b0011100100101: color_data = 12'b001110100111;
		13'b0011100101101: color_data = 12'b001110100111;
		13'b0011100101110: color_data = 12'b001110100111;
		13'b0011100110000: color_data = 12'b001110100111;
		13'b0011100111000: color_data = 12'b001110100111;
		13'b0011100111001: color_data = 12'b001110100111;
		13'b0011100111010: color_data = 12'b001110100111;
		13'b0011100111100: color_data = 12'b001110100111;
		13'b0011101000011: color_data = 12'b001110100111;
		13'b0011101000100: color_data = 12'b001110100111;
		13'b0011101000110: color_data = 12'b001110100111;
		13'b0011101001000: color_data = 12'b001110100111;
		13'b0011101001001: color_data = 12'b001110100111;
		13'b0011101001011: color_data = 12'b001110100111;
		13'b0011101001100: color_data = 12'b001110100111;
		13'b0011101001101: color_data = 12'b001110100111;
		13'b0011101010101: color_data = 12'b001110100111;
		13'b0011101010110: color_data = 12'b001110100111;
		13'b0011101011000: color_data = 12'b001110100111;
		13'b0011101011010: color_data = 12'b001110100111;
		13'b0011101011011: color_data = 12'b001110100111;
		13'b0011101011100: color_data = 12'b001110100111;
		13'b0011101100100: color_data = 12'b001110100111;
		13'b0011101100101: color_data = 12'b001110100111;
		13'b0011101100110: color_data = 12'b001110100111;
		13'b0011101101000: color_data = 12'b001110100111;
		13'b0011101101010: color_data = 12'b001110100111;
		13'b0011101101011: color_data = 12'b001110100111;
		13'b0011101101101: color_data = 12'b001110100111;
		13'b0011110000011: color_data = 12'b001110100111;
		13'b0011110000101: color_data = 12'b001110100111;
		13'b0011110000110: color_data = 12'b001110100111;
		13'b0011110000111: color_data = 12'b001110100111;
		13'b0100000000000: color_data = 12'b001110100111;
		13'b0100000000001: color_data = 12'b001110100111;
		13'b0100000000010: color_data = 12'b001110100111;
		13'b0100000000100: color_data = 12'b001110100111;
		13'b0100000010000: color_data = 12'b001110100111;
		13'b0100000010001: color_data = 12'b001110100111;
		13'b0100000010010: color_data = 12'b001110100111;
		13'b0100000011010: color_data = 12'b001110100111;
		13'b0100000011100: color_data = 12'b001110100111;
		13'b0100000011101: color_data = 12'b001110100111;
		13'b0100000011110: color_data = 12'b001110100111;
		13'b0100000100000: color_data = 12'b001110100111;
		13'b0100000100001: color_data = 12'b001110100111;
		13'b0100000100011: color_data = 12'b001110100111;
		13'b0100000100100: color_data = 12'b001110100111;
		13'b0100000100101: color_data = 12'b001110100111;
		13'b0100000100110: color_data = 12'b001110100111;
		13'b0100000101101: color_data = 12'b001110100111;
		13'b0100000101110: color_data = 12'b001110100111;
		13'b0100000110000: color_data = 12'b001110100111;
		13'b0100000111000: color_data = 12'b001110100111;
		13'b0100000111001: color_data = 12'b001110100111;
		13'b0100000111010: color_data = 12'b001110100111;
		13'b0100000111100: color_data = 12'b001110100111;
		13'b0100001000011: color_data = 12'b001110100111;
		13'b0100001000100: color_data = 12'b001110100111;
		13'b0100001000110: color_data = 12'b001110100111;
		13'b0100001001000: color_data = 12'b001110100111;
		13'b0100001001001: color_data = 12'b001110100111;
		13'b0100001001011: color_data = 12'b001110100111;
		13'b0100001001100: color_data = 12'b001110100111;
		13'b0100001001101: color_data = 12'b001110100111;
		13'b0100001001110: color_data = 12'b001110100111;
		13'b0100001010101: color_data = 12'b001110100111;
		13'b0100001010110: color_data = 12'b001110100111;
		13'b0100001011000: color_data = 12'b001110100111;
		13'b0100001011010: color_data = 12'b001110100111;
		13'b0100001011011: color_data = 12'b001110100111;
		13'b0100001011100: color_data = 12'b001110100111;
		13'b0100001100100: color_data = 12'b001110100111;
		13'b0100001100101: color_data = 12'b001110100111;
		13'b0100001100110: color_data = 12'b001110100111;
		13'b0100001101000: color_data = 12'b001110100111;
		13'b0100001101010: color_data = 12'b001110100111;
		13'b0100001101011: color_data = 12'b001110100111;
		13'b0100001101101: color_data = 12'b001110100111;
		13'b0100010000011: color_data = 12'b001110100111;
		13'b0100010000101: color_data = 12'b001110100111;
		13'b0100010000110: color_data = 12'b001110100111;
		13'b0100010000111: color_data = 12'b001110100111;
		13'b0100100000000: color_data = 12'b001110100111;
		13'b0100100000001: color_data = 12'b001110100111;
		13'b0100100000010: color_data = 12'b001110100111;
		13'b0100100000100: color_data = 12'b001110100111;
		13'b0100100010000: color_data = 12'b001110100111;
		13'b0100100010001: color_data = 12'b001110100111;
		13'b0100100010010: color_data = 12'b001110100111;
		13'b0100100011010: color_data = 12'b001110100111;
		13'b0100100011100: color_data = 12'b001110100111;
		13'b0100100011101: color_data = 12'b001110100111;
		13'b0100100011110: color_data = 12'b001110100111;
		13'b0100100100000: color_data = 12'b001110100111;
		13'b0100100100001: color_data = 12'b001110100111;
		13'b0100100100011: color_data = 12'b001110100111;
		13'b0100100100100: color_data = 12'b001110100111;
		13'b0100100100101: color_data = 12'b001110100111;
		13'b0100100100110: color_data = 12'b001110100111;
		13'b0100100101101: color_data = 12'b001110100111;
		13'b0100100101110: color_data = 12'b001110100111;
		13'b0100100110000: color_data = 12'b001110100111;
		13'b0100100111000: color_data = 12'b001110100111;
		13'b0100100111001: color_data = 12'b001110100111;
		13'b0100100111010: color_data = 12'b001110100111;
		13'b0100100111100: color_data = 12'b001110100111;
		13'b0100101000011: color_data = 12'b001110100111;
		13'b0100101000100: color_data = 12'b001110100111;
		13'b0100101000110: color_data = 12'b001110100111;
		13'b0100101001000: color_data = 12'b001110100111;
		13'b0100101001001: color_data = 12'b001110100111;
		13'b0100101001011: color_data = 12'b001110100111;
		13'b0100101001100: color_data = 12'b001110100111;
		13'b0100101001101: color_data = 12'b001110100111;
		13'b0100101001110: color_data = 12'b001110100111;
		13'b0100101010101: color_data = 12'b001110100111;
		13'b0100101010110: color_data = 12'b001110100111;
		13'b0100101011000: color_data = 12'b001110100111;
		13'b0100101011010: color_data = 12'b001110100111;
		13'b0100101011011: color_data = 12'b001110100111;
		13'b0100101011100: color_data = 12'b001110100111;
		13'b0100101100100: color_data = 12'b001110100111;
		13'b0100101100101: color_data = 12'b001110100111;
		13'b0100101100110: color_data = 12'b001110100111;
		13'b0100101101000: color_data = 12'b001110100111;
		13'b0100101101010: color_data = 12'b001110100111;
		13'b0100101101011: color_data = 12'b001110100111;
		13'b0100101101101: color_data = 12'b001110100111;
		13'b0100110000011: color_data = 12'b001110100111;
		13'b0100110000101: color_data = 12'b001110100111;
		13'b0100110000110: color_data = 12'b001110100111;
		13'b0100110000111: color_data = 12'b001110100111;
		13'b0101000000000: color_data = 12'b001110100111;
		13'b0101000000001: color_data = 12'b001110100111;
		13'b0101000000010: color_data = 12'b001110100111;
		13'b0101000000100: color_data = 12'b001110100111;
		13'b0101000010000: color_data = 12'b001110100111;
		13'b0101000010001: color_data = 12'b001110100111;
		13'b0101000010010: color_data = 12'b001110100111;
		13'b0101000011010: color_data = 12'b001110100111;
		13'b0101000011100: color_data = 12'b001110100111;
		13'b0101000011101: color_data = 12'b001110100111;
		13'b0101000011110: color_data = 12'b001110100111;
		13'b0101000100000: color_data = 12'b001110100111;
		13'b0101000100001: color_data = 12'b001110100111;
		13'b0101000100011: color_data = 12'b001110100111;
		13'b0101000100101: color_data = 12'b001110100111;
		13'b0101000100110: color_data = 12'b001110100111;
		13'b0101000100111: color_data = 12'b001110100111;
		13'b0101000101101: color_data = 12'b001110100111;
		13'b0101000101110: color_data = 12'b001110100111;
		13'b0101000110000: color_data = 12'b001110100111;
		13'b0101000111000: color_data = 12'b001110100111;
		13'b0101000111001: color_data = 12'b001110100111;
		13'b0101000111010: color_data = 12'b001110100111;
		13'b0101000111100: color_data = 12'b001110100111;
		13'b0101001000011: color_data = 12'b001110100111;
		13'b0101001000100: color_data = 12'b001110100111;
		13'b0101001000110: color_data = 12'b001110100111;
		13'b0101001001000: color_data = 12'b001110100111;
		13'b0101001001001: color_data = 12'b001110100111;
		13'b0101001001011: color_data = 12'b001110100111;
		13'b0101001001101: color_data = 12'b001110100111;
		13'b0101001001110: color_data = 12'b001110100111;
		13'b0101001001111: color_data = 12'b001110100111;
		13'b0101001010101: color_data = 12'b001110100111;
		13'b0101001010110: color_data = 12'b001110100111;
		13'b0101001011000: color_data = 12'b001110100111;
		13'b0101001011010: color_data = 12'b001110100111;
		13'b0101001011011: color_data = 12'b001110100111;
		13'b0101001011100: color_data = 12'b001110100111;
		13'b0101001100100: color_data = 12'b001110100111;
		13'b0101001100101: color_data = 12'b001110100111;
		13'b0101001100110: color_data = 12'b001110100111;
		13'b0101001101000: color_data = 12'b001110100111;
		13'b0101001101010: color_data = 12'b001110100111;
		13'b0101001101011: color_data = 12'b001110100111;
		13'b0101001101101: color_data = 12'b001110100111;
		13'b0101010000011: color_data = 12'b001110100111;
		13'b0101010000101: color_data = 12'b001110100111;
		13'b0101010000110: color_data = 12'b001110100111;
		13'b0101010000111: color_data = 12'b001110100111;
		13'b0101100000000: color_data = 12'b001110100111;
		13'b0101100000001: color_data = 12'b001110100111;
		13'b0101100000010: color_data = 12'b001110100111;
		13'b0101100000100: color_data = 12'b001110100111;
		13'b0101100010000: color_data = 12'b001110100111;
		13'b0101100010001: color_data = 12'b001110100111;
		13'b0101100010010: color_data = 12'b001110100111;
		13'b0101100011010: color_data = 12'b001110100111;
		13'b0101100011100: color_data = 12'b001110100111;
		13'b0101100011101: color_data = 12'b001110100111;
		13'b0101100011110: color_data = 12'b001110100111;
		13'b0101100100000: color_data = 12'b001110100111;
		13'b0101100100001: color_data = 12'b001110100111;
		13'b0101100100011: color_data = 12'b001110100111;
		13'b0101100100101: color_data = 12'b001110100111;
		13'b0101100100110: color_data = 12'b001110100111;
		13'b0101100100111: color_data = 12'b001110100111;
		13'b0101100101101: color_data = 12'b001110100111;
		13'b0101100101110: color_data = 12'b001110100111;
		13'b0101100110000: color_data = 12'b001110100111;
		13'b0101100111000: color_data = 12'b001110100111;
		13'b0101100111001: color_data = 12'b001110100111;
		13'b0101100111010: color_data = 12'b001110100111;
		13'b0101100111100: color_data = 12'b001110100111;
		13'b0101101000011: color_data = 12'b001110100111;
		13'b0101101000100: color_data = 12'b001110100111;
		13'b0101101000110: color_data = 12'b001110100111;
		13'b0101101001000: color_data = 12'b001110100111;
		13'b0101101001001: color_data = 12'b001110100111;
		13'b0101101001011: color_data = 12'b001110100111;
		13'b0101101001101: color_data = 12'b001110100111;
		13'b0101101001110: color_data = 12'b001110100111;
		13'b0101101001111: color_data = 12'b001110100111;
		13'b0101101010101: color_data = 12'b001110100111;
		13'b0101101010110: color_data = 12'b001110100111;
		13'b0101101011000: color_data = 12'b001110100111;
		13'b0101101011010: color_data = 12'b001110100111;
		13'b0101101011011: color_data = 12'b001110100111;
		13'b0101101011100: color_data = 12'b001110100111;
		13'b0101101100100: color_data = 12'b001110100111;
		13'b0101101100101: color_data = 12'b001110100111;
		13'b0101101100110: color_data = 12'b001110100111;
		13'b0101101101000: color_data = 12'b001110100111;
		13'b0101101101010: color_data = 12'b001110100111;
		13'b0101101101011: color_data = 12'b001110100111;
		13'b0101101101100: color_data = 12'b001110100111;
		13'b0101101101101: color_data = 12'b001110100111;
		13'b0101101101110: color_data = 12'b001110100111;
		13'b0101101101111: color_data = 12'b001110100111;
		13'b0101101110000: color_data = 12'b001110100111;
		13'b0101101110001: color_data = 12'b001110100111;
		13'b0101101110010: color_data = 12'b001110100111;
		13'b0101101110011: color_data = 12'b001110100111;
		13'b0101101110100: color_data = 12'b001110100111;
		13'b0101101110101: color_data = 12'b001110100111;
		13'b0101110000011: color_data = 12'b001110100111;
		13'b0101110000100: color_data = 12'b001110100111;
		13'b0101110000101: color_data = 12'b001110100111;
		13'b0101110000110: color_data = 12'b001110100111;
		13'b0110000000000: color_data = 12'b001110100111;
		13'b0110000000001: color_data = 12'b001110100111;
		13'b0110000000010: color_data = 12'b001110100111;
		13'b0110000000100: color_data = 12'b001110100111;
		13'b0110000010000: color_data = 12'b001110100111;
		13'b0110000010001: color_data = 12'b001110100111;
		13'b0110000010010: color_data = 12'b001110100111;
		13'b0110000011010: color_data = 12'b001110100111;
		13'b0110000011100: color_data = 12'b001110100111;
		13'b0110000011101: color_data = 12'b001110100111;
		13'b0110000011110: color_data = 12'b001110100111;
		13'b0110000100000: color_data = 12'b001110100111;
		13'b0110000100001: color_data = 12'b001110100111;
		13'b0110000100011: color_data = 12'b001110100111;
		13'b0110000100110: color_data = 12'b001110100111;
		13'b0110000100111: color_data = 12'b001110100111;
		13'b0110000101000: color_data = 12'b001110100111;
		13'b0110000101101: color_data = 12'b001110100111;
		13'b0110000101110: color_data = 12'b001110100111;
		13'b0110000110000: color_data = 12'b001110100111;
		13'b0110000111000: color_data = 12'b001110100111;
		13'b0110000111001: color_data = 12'b001110100111;
		13'b0110000111010: color_data = 12'b001110100111;
		13'b0110000111100: color_data = 12'b001110100111;
		13'b0110001000011: color_data = 12'b001110100111;
		13'b0110001000100: color_data = 12'b001110100111;
		13'b0110001000110: color_data = 12'b001110100111;
		13'b0110001001000: color_data = 12'b001110100111;
		13'b0110001001001: color_data = 12'b001110100111;
		13'b0110001001011: color_data = 12'b001110100111;
		13'b0110001001110: color_data = 12'b001110100111;
		13'b0110001001111: color_data = 12'b001110100111;
		13'b0110001010000: color_data = 12'b001110100111;
		13'b0110001010101: color_data = 12'b001110100111;
		13'b0110001010110: color_data = 12'b001110100111;
		13'b0110001011000: color_data = 12'b001110100111;
		13'b0110001011010: color_data = 12'b001110100111;
		13'b0110001011011: color_data = 12'b001110100111;
		13'b0110001011100: color_data = 12'b001110100111;
		13'b0110001100100: color_data = 12'b001110100111;
		13'b0110001100101: color_data = 12'b001110100111;
		13'b0110001100110: color_data = 12'b001110100111;
		13'b0110001101000: color_data = 12'b001110100111;
		13'b0110001101010: color_data = 12'b001110100111;
		13'b0110001101011: color_data = 12'b001110100111;
		13'b0110001101100: color_data = 12'b001110100111;
		13'b0110001101101: color_data = 12'b001110100111;
		13'b0110001101110: color_data = 12'b001110100111;
		13'b0110001101111: color_data = 12'b001110100111;
		13'b0110001110000: color_data = 12'b001110100111;
		13'b0110001110001: color_data = 12'b001110100111;
		13'b0110001110010: color_data = 12'b001110100111;
		13'b0110001110011: color_data = 12'b001110100111;
		13'b0110001110100: color_data = 12'b001110100111;
		13'b0110001110101: color_data = 12'b001110100111;
		13'b0110010000011: color_data = 12'b001110100111;
		13'b0110010000100: color_data = 12'b001110100111;
		13'b0110010000101: color_data = 12'b001110100111;
		13'b0110100000000: color_data = 12'b001110100111;
		13'b0110100000001: color_data = 12'b001110100111;
		13'b0110100000010: color_data = 12'b001110100111;
		13'b0110100000100: color_data = 12'b001110100111;
		13'b0110100010000: color_data = 12'b001110100111;
		13'b0110100010001: color_data = 12'b001110100111;
		13'b0110100010010: color_data = 12'b001110100111;
		13'b0110100011010: color_data = 12'b001110100111;
		13'b0110100011100: color_data = 12'b001110100111;
		13'b0110100011101: color_data = 12'b001110100111;
		13'b0110100011110: color_data = 12'b001110100111;
		13'b0110100100000: color_data = 12'b001110100111;
		13'b0110100100001: color_data = 12'b001110100111;
		13'b0110100100011: color_data = 12'b001110100111;
		13'b0110100100110: color_data = 12'b001110100111;
		13'b0110100100111: color_data = 12'b001110100111;
		13'b0110100101000: color_data = 12'b001110100111;
		13'b0110100101101: color_data = 12'b001110100111;
		13'b0110100101110: color_data = 12'b001110100111;
		13'b0110100110000: color_data = 12'b001110100111;
		13'b0110100111000: color_data = 12'b001110100111;
		13'b0110100111001: color_data = 12'b001110100111;
		13'b0110100111010: color_data = 12'b001110100111;
		13'b0110100111100: color_data = 12'b001110100111;
		13'b0110101000011: color_data = 12'b001110100111;
		13'b0110101000100: color_data = 12'b001110100111;
		13'b0110101000110: color_data = 12'b001110100111;
		13'b0110101001000: color_data = 12'b001110100111;
		13'b0110101001001: color_data = 12'b001110100111;
		13'b0110101001011: color_data = 12'b001110100111;
		13'b0110101001110: color_data = 12'b001110100111;
		13'b0110101001111: color_data = 12'b001110100111;
		13'b0110101010000: color_data = 12'b001110100111;
		13'b0110101010101: color_data = 12'b001110100111;
		13'b0110101010110: color_data = 12'b001110100111;
		13'b0110101011000: color_data = 12'b001110100111;
		13'b0110101011010: color_data = 12'b001110100111;
		13'b0110101011011: color_data = 12'b001110100111;
		13'b0110101011100: color_data = 12'b001110100111;
		13'b0110101100100: color_data = 12'b001110100111;
		13'b0110101100101: color_data = 12'b001110100111;
		13'b0110101100110: color_data = 12'b001110100111;
		13'b0110101101000: color_data = 12'b001110100111;
		13'b0110101101010: color_data = 12'b001110100111;
		13'b0110101101011: color_data = 12'b001110100111;
		13'b0110101101100: color_data = 12'b001110100111;
		13'b0110101101101: color_data = 12'b001110100111;
		13'b0110101101110: color_data = 12'b001110100111;
		13'b0110101101111: color_data = 12'b001110100111;
		13'b0110101110000: color_data = 12'b001110100111;
		13'b0110101110001: color_data = 12'b001110100111;
		13'b0110101110010: color_data = 12'b001110100111;
		13'b0110101110011: color_data = 12'b001110100111;
		13'b0110101110100: color_data = 12'b001110100111;
		13'b0110101110101: color_data = 12'b001110100111;
		13'b0110110000010: color_data = 12'b001110100111;
		13'b0110110000011: color_data = 12'b001110100111;
		13'b0110110000100: color_data = 12'b001110100111;
		13'b0111000000000: color_data = 12'b001110100111;
		13'b0111000000001: color_data = 12'b001110100111;
		13'b0111000000010: color_data = 12'b001110100111;
		13'b0111000000100: color_data = 12'b001110100111;
		13'b0111000010000: color_data = 12'b001110100111;
		13'b0111000010001: color_data = 12'b001110100111;
		13'b0111000010010: color_data = 12'b001110100111;
		13'b0111000011010: color_data = 12'b001110100111;
		13'b0111000011100: color_data = 12'b001110100111;
		13'b0111000011101: color_data = 12'b001110100111;
		13'b0111000011110: color_data = 12'b001110100111;
		13'b0111000100000: color_data = 12'b001110100111;
		13'b0111000100001: color_data = 12'b001110100111;
		13'b0111000100011: color_data = 12'b001110100111;
		13'b0111000100111: color_data = 12'b001110100111;
		13'b0111000101000: color_data = 12'b001110100111;
		13'b0111000101001: color_data = 12'b001110100111;
		13'b0111000101101: color_data = 12'b001110100111;
		13'b0111000101110: color_data = 12'b001110100111;
		13'b0111000110000: color_data = 12'b001110100111;
		13'b0111000111000: color_data = 12'b001110100111;
		13'b0111000111001: color_data = 12'b001110100111;
		13'b0111000111010: color_data = 12'b001110100111;
		13'b0111000111100: color_data = 12'b001110100111;
		13'b0111001000011: color_data = 12'b001110100111;
		13'b0111001000100: color_data = 12'b001110100111;
		13'b0111001000110: color_data = 12'b001110100111;
		13'b0111001001000: color_data = 12'b001110100111;
		13'b0111001001001: color_data = 12'b001110100111;
		13'b0111001001011: color_data = 12'b001110100111;
		13'b0111001001111: color_data = 12'b001110100111;
		13'b0111001010000: color_data = 12'b001110100111;
		13'b0111001010001: color_data = 12'b001110100111;
		13'b0111001010101: color_data = 12'b001110100111;
		13'b0111001010110: color_data = 12'b001110100111;
		13'b0111001011000: color_data = 12'b001110100111;
		13'b0111001011010: color_data = 12'b001110100111;
		13'b0111001011011: color_data = 12'b001110100111;
		13'b0111001011100: color_data = 12'b001110100111;
		13'b0111001100100: color_data = 12'b001110100111;
		13'b0111001100101: color_data = 12'b001110100111;
		13'b0111001100110: color_data = 12'b001110100111;
		13'b0111001101000: color_data = 12'b001110100111;
		13'b0111001101010: color_data = 12'b001110100111;
		13'b0111001101011: color_data = 12'b001110100111;
		13'b0111001101101: color_data = 12'b001110100111;
		13'b0111010000001: color_data = 12'b001110100111;
		13'b0111010000010: color_data = 12'b001110100111;
		13'b0111010000011: color_data = 12'b001110100111;
		13'b0111100000000: color_data = 12'b001110100111;
		13'b0111100000001: color_data = 12'b001110100111;
		13'b0111100000010: color_data = 12'b001110100111;
		13'b0111100000100: color_data = 12'b001110100111;
		13'b0111100010000: color_data = 12'b001110100111;
		13'b0111100010001: color_data = 12'b001110100111;
		13'b0111100010010: color_data = 12'b001110100111;
		13'b0111100011010: color_data = 12'b001110100111;
		13'b0111100011100: color_data = 12'b001110100111;
		13'b0111100011101: color_data = 12'b001110100111;
		13'b0111100011110: color_data = 12'b001110100111;
		13'b0111100100000: color_data = 12'b001110100111;
		13'b0111100100001: color_data = 12'b001110100111;
		13'b0111100100011: color_data = 12'b001110100111;
		13'b0111100100111: color_data = 12'b001110100111;
		13'b0111100101000: color_data = 12'b001110100111;
		13'b0111100101001: color_data = 12'b001110100111;
		13'b0111100101101: color_data = 12'b001110100111;
		13'b0111100101110: color_data = 12'b001110100111;
		13'b0111100110000: color_data = 12'b001110100111;
		13'b0111100111000: color_data = 12'b001110100111;
		13'b0111100111001: color_data = 12'b001110100111;
		13'b0111100111010: color_data = 12'b001110100111;
		13'b0111100111100: color_data = 12'b001110100111;
		13'b0111101000011: color_data = 12'b001110100111;
		13'b0111101000100: color_data = 12'b001110100111;
		13'b0111101000110: color_data = 12'b001110100111;
		13'b0111101001000: color_data = 12'b001110100111;
		13'b0111101001001: color_data = 12'b001110100111;
		13'b0111101001011: color_data = 12'b001110100111;
		13'b0111101001111: color_data = 12'b001110100111;
		13'b0111101010000: color_data = 12'b001110100111;
		13'b0111101010001: color_data = 12'b001110100111;
		13'b0111101010101: color_data = 12'b001110100111;
		13'b0111101010110: color_data = 12'b001110100111;
		13'b0111101011000: color_data = 12'b001110100111;
		13'b0111101011010: color_data = 12'b001110100111;
		13'b0111101011011: color_data = 12'b001110100111;
		13'b0111101011100: color_data = 12'b001110100111;
		13'b0111101100100: color_data = 12'b001110100111;
		13'b0111101100101: color_data = 12'b001110100111;
		13'b0111101100110: color_data = 12'b001110100111;
		13'b0111101101000: color_data = 12'b001110100111;
		13'b0111101101010: color_data = 12'b001110100111;
		13'b0111101101011: color_data = 12'b001110100111;
		13'b0111101101101: color_data = 12'b001110100111;
		13'b0111110000000: color_data = 12'b001110100111;
		13'b0111110000001: color_data = 12'b001110100111;
		13'b0111110000010: color_data = 12'b001110100111;
		13'b1000000000000: color_data = 12'b001110100111;
		13'b1000000000001: color_data = 12'b001110100111;
		13'b1000000000010: color_data = 12'b001110100111;
		13'b1000000000100: color_data = 12'b001110100111;
		13'b1000000010000: color_data = 12'b001110100111;
		13'b1000000010001: color_data = 12'b001110100111;
		13'b1000000010010: color_data = 12'b001110100111;
		13'b1000000011010: color_data = 12'b001110100111;
		13'b1000000011100: color_data = 12'b001110100111;
		13'b1000000011101: color_data = 12'b001110100111;
		13'b1000000011110: color_data = 12'b001110100111;
		13'b1000000100000: color_data = 12'b001110100111;
		13'b1000000100001: color_data = 12'b001110100111;
		13'b1000000100011: color_data = 12'b001110100111;
		13'b1000000101000: color_data = 12'b001110100111;
		13'b1000000101001: color_data = 12'b001110100111;
		13'b1000000101010: color_data = 12'b001110100111;
		13'b1000000101101: color_data = 12'b001110100111;
		13'b1000000101110: color_data = 12'b001110100111;
		13'b1000000110000: color_data = 12'b001110100111;
		13'b1000000111000: color_data = 12'b001110100111;
		13'b1000000111001: color_data = 12'b001110100111;
		13'b1000000111010: color_data = 12'b001110100111;
		13'b1000000111100: color_data = 12'b001110100111;
		13'b1000001000011: color_data = 12'b001110100111;
		13'b1000001000100: color_data = 12'b001110100111;
		13'b1000001000110: color_data = 12'b001110100111;
		13'b1000001001000: color_data = 12'b001110100111;
		13'b1000001001001: color_data = 12'b001110100111;
		13'b1000001001011: color_data = 12'b001110100111;
		13'b1000001010000: color_data = 12'b001110100111;
		13'b1000001010001: color_data = 12'b001110100111;
		13'b1000001010010: color_data = 12'b001110100111;
		13'b1000001010101: color_data = 12'b001110100111;
		13'b1000001010110: color_data = 12'b001110100111;
		13'b1000001011000: color_data = 12'b001110100111;
		13'b1000001011010: color_data = 12'b001110100111;
		13'b1000001011011: color_data = 12'b001110100111;
		13'b1000001011100: color_data = 12'b001110100111;
		13'b1000001100100: color_data = 12'b001110100111;
		13'b1000001100101: color_data = 12'b001110100111;
		13'b1000001100110: color_data = 12'b001110100111;
		13'b1000001101000: color_data = 12'b001110100111;
		13'b1000001101010: color_data = 12'b001110100111;
		13'b1000001101011: color_data = 12'b001110100111;
		13'b1000001101101: color_data = 12'b001110100111;
		13'b1000010000000: color_data = 12'b001110100111;
		13'b1000010000001: color_data = 12'b001110100111;
		13'b1000010000010: color_data = 12'b001110100111;
		13'b1000100000000: color_data = 12'b001110100111;
		13'b1000100000001: color_data = 12'b001110100111;
		13'b1000100000010: color_data = 12'b001110100111;
		13'b1000100000100: color_data = 12'b001110100111;
		13'b1000100010000: color_data = 12'b001110100111;
		13'b1000100010001: color_data = 12'b001110100111;
		13'b1000100010010: color_data = 12'b001110100111;
		13'b1000100011010: color_data = 12'b001110100111;
		13'b1000100011100: color_data = 12'b001110100111;
		13'b1000100011101: color_data = 12'b001110100111;
		13'b1000100011110: color_data = 12'b001110100111;
		13'b1000100100000: color_data = 12'b001110100111;
		13'b1000100100001: color_data = 12'b001110100111;
		13'b1000100100011: color_data = 12'b001110100111;
		13'b1000100101000: color_data = 12'b001110100111;
		13'b1000100101001: color_data = 12'b001110100111;
		13'b1000100101010: color_data = 12'b001110100111;
		13'b1000100101101: color_data = 12'b001110100111;
		13'b1000100101110: color_data = 12'b001110100111;
		13'b1000100110000: color_data = 12'b001110100111;
		13'b1000100111000: color_data = 12'b001110100111;
		13'b1000100111001: color_data = 12'b001110100111;
		13'b1000100111010: color_data = 12'b001110100111;
		13'b1000100111100: color_data = 12'b001110100111;
		13'b1000101000011: color_data = 12'b001110100111;
		13'b1000101000100: color_data = 12'b001110100111;
		13'b1000101000110: color_data = 12'b001110100111;
		13'b1000101001000: color_data = 12'b001110100111;
		13'b1000101001001: color_data = 12'b001110100111;
		13'b1000101001011: color_data = 12'b001110100111;
		13'b1000101010000: color_data = 12'b001110100111;
		13'b1000101010001: color_data = 12'b001110100111;
		13'b1000101010010: color_data = 12'b001110100111;
		13'b1000101010101: color_data = 12'b001110100111;
		13'b1000101010110: color_data = 12'b001110100111;
		13'b1000101011000: color_data = 12'b001110100111;
		13'b1000101011010: color_data = 12'b001110100111;
		13'b1000101011011: color_data = 12'b001110100111;
		13'b1000101011100: color_data = 12'b001110100111;
		13'b1000101100100: color_data = 12'b001110100111;
		13'b1000101100101: color_data = 12'b001110100111;
		13'b1000101100110: color_data = 12'b001110100111;
		13'b1000101101000: color_data = 12'b001110100111;
		13'b1000101101010: color_data = 12'b001110100111;
		13'b1000101101011: color_data = 12'b001110100111;
		13'b1000101101101: color_data = 12'b001110100111;
		13'b1000110000000: color_data = 12'b001110100111;
		13'b1000110000001: color_data = 12'b001110100111;
		13'b1000110000010: color_data = 12'b001110100111;
		13'b1001000000000: color_data = 12'b001110100111;
		13'b1001000000001: color_data = 12'b001110100111;
		13'b1001000000010: color_data = 12'b001110100111;
		13'b1001000000100: color_data = 12'b001110100111;
		13'b1001000001100: color_data = 12'b001110100111;
		13'b1001000001101: color_data = 12'b001110100111;
		13'b1001000001110: color_data = 12'b001110100111;
		13'b1001000010000: color_data = 12'b001110100111;
		13'b1001000010001: color_data = 12'b001110100111;
		13'b1001000010010: color_data = 12'b001110100111;
		13'b1001000011010: color_data = 12'b001110100111;
		13'b1001000011100: color_data = 12'b001110100111;
		13'b1001000011101: color_data = 12'b001110100111;
		13'b1001000011110: color_data = 12'b001110100111;
		13'b1001000100000: color_data = 12'b001110100111;
		13'b1001000100001: color_data = 12'b001110100111;
		13'b1001000100011: color_data = 12'b001110100111;
		13'b1001000101001: color_data = 12'b001110100111;
		13'b1001000101010: color_data = 12'b001110100111;
		13'b1001000101011: color_data = 12'b001110100111;
		13'b1001000101101: color_data = 12'b001110100111;
		13'b1001000101110: color_data = 12'b001110100111;
		13'b1001000110000: color_data = 12'b001110100111;
		13'b1001000111000: color_data = 12'b001110100111;
		13'b1001000111001: color_data = 12'b001110100111;
		13'b1001000111010: color_data = 12'b001110100111;
		13'b1001000111100: color_data = 12'b001110100111;
		13'b1001001000011: color_data = 12'b001110100111;
		13'b1001001000100: color_data = 12'b001110100111;
		13'b1001001000110: color_data = 12'b001110100111;
		13'b1001001001000: color_data = 12'b001110100111;
		13'b1001001001001: color_data = 12'b001110100111;
		13'b1001001001011: color_data = 12'b001110100111;
		13'b1001001010001: color_data = 12'b001110100111;
		13'b1001001010010: color_data = 12'b001110100111;
		13'b1001001010011: color_data = 12'b001110100111;
		13'b1001001010101: color_data = 12'b001110100111;
		13'b1001001010110: color_data = 12'b001110100111;
		13'b1001001011000: color_data = 12'b001110100111;
		13'b1001001011010: color_data = 12'b001110100111;
		13'b1001001011011: color_data = 12'b001110100111;
		13'b1001001011100: color_data = 12'b001110100111;
		13'b1001001100100: color_data = 12'b001110100111;
		13'b1001001100101: color_data = 12'b001110100111;
		13'b1001001100110: color_data = 12'b001110100111;
		13'b1001001101000: color_data = 12'b001110100111;
		13'b1001001101010: color_data = 12'b001110100111;
		13'b1001001101011: color_data = 12'b001110100111;
		13'b1001001101101: color_data = 12'b001110100111;
		13'b1001010000000: color_data = 12'b001110100111;
		13'b1001010000001: color_data = 12'b001110100111;
		13'b1001010000010: color_data = 12'b001110100111;
		13'b1001100000000: color_data = 12'b001110100111;
		13'b1001100000001: color_data = 12'b001110100111;
		13'b1001100000010: color_data = 12'b001110100111;
		13'b1001100000100: color_data = 12'b001110100111;
		13'b1001100001100: color_data = 12'b001110100111;
		13'b1001100001101: color_data = 12'b001110100111;
		13'b1001100001110: color_data = 12'b001110100111;
		13'b1001100010000: color_data = 12'b001110100111;
		13'b1001100010001: color_data = 12'b001110100111;
		13'b1001100010010: color_data = 12'b001110100111;
		13'b1001100011010: color_data = 12'b001110100111;
		13'b1001100011100: color_data = 12'b001110100111;
		13'b1001100011101: color_data = 12'b001110100111;
		13'b1001100011110: color_data = 12'b001110100111;
		13'b1001100100000: color_data = 12'b001110100111;
		13'b1001100100001: color_data = 12'b001110100111;
		13'b1001100100011: color_data = 12'b001110100111;
		13'b1001100101001: color_data = 12'b001110100111;
		13'b1001100101010: color_data = 12'b001110100111;
		13'b1001100101011: color_data = 12'b001110100111;
		13'b1001100101101: color_data = 12'b001110100111;
		13'b1001100101110: color_data = 12'b001110100111;
		13'b1001100110000: color_data = 12'b001110100111;
		13'b1001100111000: color_data = 12'b001110100111;
		13'b1001100111001: color_data = 12'b001110100111;
		13'b1001100111010: color_data = 12'b001110100111;
		13'b1001100111100: color_data = 12'b001110100111;
		13'b1001101000011: color_data = 12'b001110100111;
		13'b1001101000100: color_data = 12'b001110100111;
		13'b1001101000110: color_data = 12'b001110100111;
		13'b1001101001000: color_data = 12'b001110100111;
		13'b1001101001001: color_data = 12'b001110100111;
		13'b1001101001011: color_data = 12'b001110100111;
		13'b1001101010001: color_data = 12'b001110100111;
		13'b1001101010010: color_data = 12'b001110100111;
		13'b1001101010011: color_data = 12'b001110100111;
		13'b1001101010101: color_data = 12'b001110100111;
		13'b1001101010110: color_data = 12'b001110100111;
		13'b1001101011000: color_data = 12'b001110100111;
		13'b1001101011010: color_data = 12'b001110100111;
		13'b1001101011011: color_data = 12'b001110100111;
		13'b1001101011100: color_data = 12'b001110100111;
		13'b1001101100100: color_data = 12'b001110100111;
		13'b1001101100101: color_data = 12'b001110100111;
		13'b1001101100110: color_data = 12'b001110100111;
		13'b1001101101000: color_data = 12'b001110100111;
		13'b1001101101010: color_data = 12'b001110100111;
		13'b1001101101011: color_data = 12'b001110100111;
		13'b1001101101101: color_data = 12'b001110100111;
		13'b1010000000001: color_data = 12'b001110100111;
		13'b1010000000010: color_data = 12'b001110100111;
		13'b1010000000011: color_data = 12'b001110100111;
		13'b1010000000100: color_data = 12'b001110100111;
		13'b1010000001011: color_data = 12'b001110100111;
		13'b1010000001100: color_data = 12'b001110100111;
		13'b1010000001101: color_data = 12'b001110100111;
		13'b1010000010000: color_data = 12'b001110100111;
		13'b1010000010001: color_data = 12'b001110100111;
		13'b1010000010010: color_data = 12'b001110100111;
		13'b1010000011010: color_data = 12'b001110100111;
		13'b1010000011100: color_data = 12'b001110100111;
		13'b1010000011101: color_data = 12'b001110100111;
		13'b1010000011110: color_data = 12'b001110100111;
		13'b1010000100000: color_data = 12'b001110100111;
		13'b1010000100001: color_data = 12'b001110100111;
		13'b1010000100011: color_data = 12'b001110100111;
		13'b1010000101010: color_data = 12'b001110100111;
		13'b1010000101011: color_data = 12'b001110100111;
		13'b1010000101100: color_data = 12'b001110100111;
		13'b1010000101101: color_data = 12'b001110100111;
		13'b1010000101110: color_data = 12'b001110100111;
		13'b1010000110000: color_data = 12'b001110100111;
		13'b1010000111000: color_data = 12'b001110100111;
		13'b1010000111001: color_data = 12'b001110100111;
		13'b1010000111010: color_data = 12'b001110100111;
		13'b1010000111100: color_data = 12'b001110100111;
		13'b1010001000011: color_data = 12'b001110100111;
		13'b1010001000100: color_data = 12'b001110100111;
		13'b1010001000110: color_data = 12'b001110100111;
		13'b1010001001000: color_data = 12'b001110100111;
		13'b1010001001001: color_data = 12'b001110100111;
		13'b1010001001011: color_data = 12'b001110100111;
		13'b1010001010010: color_data = 12'b001110100111;
		13'b1010001010011: color_data = 12'b001110100111;
		13'b1010001010100: color_data = 12'b001110100111;
		13'b1010001010101: color_data = 12'b001110100111;
		13'b1010001010110: color_data = 12'b001110100111;
		13'b1010001011000: color_data = 12'b001110100111;
		13'b1010001011010: color_data = 12'b001110100111;
		13'b1010001011011: color_data = 12'b001110100111;
		13'b1010001011100: color_data = 12'b001110100111;
		13'b1010001011101: color_data = 12'b001110100111;
		13'b1010001100011: color_data = 12'b001110100111;
		13'b1010001100100: color_data = 12'b001110100111;
		13'b1010001100101: color_data = 12'b001110100111;
		13'b1010001100110: color_data = 12'b001110100111;
		13'b1010001101000: color_data = 12'b001110100111;
		13'b1010001101010: color_data = 12'b001110100111;
		13'b1010001101011: color_data = 12'b001110100111;
		13'b1010001101101: color_data = 12'b001110100111;
		13'b1010001110101: color_data = 12'b001110100111;
		13'b1010001110110: color_data = 12'b001110100111;
		13'b1010001110111: color_data = 12'b001110100111;
		13'b1010001111111: color_data = 12'b001110100111;
		13'b1010010000000: color_data = 12'b001110100111;
		13'b1010010000001: color_data = 12'b001110100111;
		13'b1010010000010: color_data = 12'b001110100111;
		13'b1010010000011: color_data = 12'b001110100111;
		13'b1010100000001: color_data = 12'b001110100111;
		13'b1010100000010: color_data = 12'b001110100111;
		13'b1010100000011: color_data = 12'b001110100111;
		13'b1010100000100: color_data = 12'b001110100111;
		13'b1010100001010: color_data = 12'b001110100111;
		13'b1010100001011: color_data = 12'b001110100111;
		13'b1010100001100: color_data = 12'b001110100111;
		13'b1010100001101: color_data = 12'b001110100111;
		13'b1010100010001: color_data = 12'b001110100111;
		13'b1010100010010: color_data = 12'b001110100111;
		13'b1010100010011: color_data = 12'b001110100111;
		13'b1010100011010: color_data = 12'b001110100111;
		13'b1010100011011: color_data = 12'b001110100111;
		13'b1010100011100: color_data = 12'b001110100111;
		13'b1010100011101: color_data = 12'b001110100111;
		13'b1010100100000: color_data = 12'b001110100111;
		13'b1010100100001: color_data = 12'b001110100111;
		13'b1010100100011: color_data = 12'b001110100111;
		13'b1010100101010: color_data = 12'b001110100111;
		13'b1010100101011: color_data = 12'b001110100111;
		13'b1010100101100: color_data = 12'b001110100111;
		13'b1010100101101: color_data = 12'b001110100111;
		13'b1010100101110: color_data = 12'b001110100111;
		13'b1010100110000: color_data = 12'b001110100111;
		13'b1010100111000: color_data = 12'b001110100111;
		13'b1010100111001: color_data = 12'b001110100111;
		13'b1010100111010: color_data = 12'b001110100111;
		13'b1010100111100: color_data = 12'b001110100111;
		13'b1010101000011: color_data = 12'b001110100111;
		13'b1010101000100: color_data = 12'b001110100111;
		13'b1010101000110: color_data = 12'b001110100111;
		13'b1010101001000: color_data = 12'b001110100111;
		13'b1010101001001: color_data = 12'b001110100111;
		13'b1010101001011: color_data = 12'b001110100111;
		13'b1010101010010: color_data = 12'b001110100111;
		13'b1010101010011: color_data = 12'b001110100111;
		13'b1010101010100: color_data = 12'b001110100111;
		13'b1010101010101: color_data = 12'b001110100111;
		13'b1010101010110: color_data = 12'b001110100111;
		13'b1010101011000: color_data = 12'b001110100111;
		13'b1010101011011: color_data = 12'b001110100111;
		13'b1010101011100: color_data = 12'b001110100111;
		13'b1010101011101: color_data = 12'b001110100111;
		13'b1010101011110: color_data = 12'b001110100111;
		13'b1010101011111: color_data = 12'b001110100111;
		13'b1010101100000: color_data = 12'b001110100111;
		13'b1010101100001: color_data = 12'b001110100111;
		13'b1010101100010: color_data = 12'b001110100111;
		13'b1010101100011: color_data = 12'b001110100111;
		13'b1010101100100: color_data = 12'b001110100111;
		13'b1010101100101: color_data = 12'b001110100111;
		13'b1010101100111: color_data = 12'b001110100111;
		13'b1010101101010: color_data = 12'b001110100111;
		13'b1010101101011: color_data = 12'b001110100111;
		13'b1010101101101: color_data = 12'b001110100111;
		13'b1010101110100: color_data = 12'b001110100111;
		13'b1010101110101: color_data = 12'b001110100111;
		13'b1010101110110: color_data = 12'b001110100111;
		13'b1010101110111: color_data = 12'b001110100111;
		13'b1010101111111: color_data = 12'b001110100111;
		13'b1010110000000: color_data = 12'b001110100111;
		13'b1010110000001: color_data = 12'b001110100111;
		13'b1010110000011: color_data = 12'b001110100111;
		13'b1011000000010: color_data = 12'b001110100111;
		13'b1011000000011: color_data = 12'b001110100111;
		13'b1011000000100: color_data = 12'b001110100111;
		13'b1011000000101: color_data = 12'b001110100111;
		13'b1011000000110: color_data = 12'b001110100111;
		13'b1011000000111: color_data = 12'b001110100111;
		13'b1011000001000: color_data = 12'b001110100111;
		13'b1011000001001: color_data = 12'b001110100111;
		13'b1011000001010: color_data = 12'b001110100111;
		13'b1011000001011: color_data = 12'b001110100111;
		13'b1011000001100: color_data = 12'b001110100111;
		13'b1011000010010: color_data = 12'b001110100111;
		13'b1011000010011: color_data = 12'b001110100111;
		13'b1011000010100: color_data = 12'b001110100111;
		13'b1011000010101: color_data = 12'b001110100111;
		13'b1011000010110: color_data = 12'b001110100111;
		13'b1011000010111: color_data = 12'b001110100111;
		13'b1011000011000: color_data = 12'b001110100111;
		13'b1011000011001: color_data = 12'b001110100111;
		13'b1011000011010: color_data = 12'b001110100111;
		13'b1011000011011: color_data = 12'b001110100111;
		13'b1011000011100: color_data = 12'b001110100111;
		13'b1011000100000: color_data = 12'b001110100111;
		13'b1011000100001: color_data = 12'b001110100111;
		13'b1011000100010: color_data = 12'b001110100111;
		13'b1011000100011: color_data = 12'b001110100111;
		13'b1011000101011: color_data = 12'b001110100111;
		13'b1011000101100: color_data = 12'b001110100111;
		13'b1011000101101: color_data = 12'b001110100111;
		13'b1011000101110: color_data = 12'b001110100111;
		13'b1011000101111: color_data = 12'b001110100111;
		13'b1011000110000: color_data = 12'b001110100111;
		13'b1011000110110: color_data = 12'b001110100111;
		13'b1011000110111: color_data = 12'b001110100111;
		13'b1011000111000: color_data = 12'b001110100111;
		13'b1011000111001: color_data = 12'b001110100111;
		13'b1011000111010: color_data = 12'b001110100111;
		13'b1011000111011: color_data = 12'b001110100111;
		13'b1011000111100: color_data = 12'b001110100111;
		13'b1011000111101: color_data = 12'b001110100111;
		13'b1011001000011: color_data = 12'b001110100111;
		13'b1011001000100: color_data = 12'b001110100111;
		13'b1011001000101: color_data = 12'b001110100111;
		13'b1011001000110: color_data = 12'b001110100111;
		13'b1011001001000: color_data = 12'b001110100111;
		13'b1011001001001: color_data = 12'b001110100111;
		13'b1011001001010: color_data = 12'b001110100111;
		13'b1011001001011: color_data = 12'b001110100111;
		13'b1011001010011: color_data = 12'b001110100111;
		13'b1011001010100: color_data = 12'b001110100111;
		13'b1011001010101: color_data = 12'b001110100111;
		13'b1011001010110: color_data = 12'b001110100111;
		13'b1011001010111: color_data = 12'b001110100111;
		13'b1011001011000: color_data = 12'b001110100111;
		13'b1011001011100: color_data = 12'b001110100111;
		13'b1011001011101: color_data = 12'b001110100111;
		13'b1011001011110: color_data = 12'b001110100111;
		13'b1011001011111: color_data = 12'b001110100111;
		13'b1011001100000: color_data = 12'b001110100111;
		13'b1011001100001: color_data = 12'b001110100111;
		13'b1011001100010: color_data = 12'b001110100111;
		13'b1011001100011: color_data = 12'b001110100111;
		13'b1011001100100: color_data = 12'b001110100111;
		13'b1011001100110: color_data = 12'b001110100111;
		13'b1011001101010: color_data = 12'b001110100111;
		13'b1011001101011: color_data = 12'b001110100111;
		13'b1011001101100: color_data = 12'b001110100111;
		13'b1011001101101: color_data = 12'b001110100111;
		13'b1011001101110: color_data = 12'b001110100111;
		13'b1011001101111: color_data = 12'b001110100111;
		13'b1011001110000: color_data = 12'b001110100111;
		13'b1011001110001: color_data = 12'b001110100111;
		13'b1011001110010: color_data = 12'b001110100111;
		13'b1011001110011: color_data = 12'b001110100111;
		13'b1011001110100: color_data = 12'b001110100111;
		13'b1011001110101: color_data = 12'b001110100111;
		13'b1011001110110: color_data = 12'b001110100111;
		13'b1011001111111: color_data = 12'b001110100111;
		13'b1011010000000: color_data = 12'b001110100111;
		13'b1011010000001: color_data = 12'b001110100111;
		13'b1011010000011: color_data = 12'b001110100111;
		13'b1011100000011: color_data = 12'b001110100111;
		13'b1011100000100: color_data = 12'b001110100111;
		13'b1011100000101: color_data = 12'b001110100111;
		13'b1011100000110: color_data = 12'b001110100111;
		13'b1011100000111: color_data = 12'b001110100111;
		13'b1011100001000: color_data = 12'b001110100111;
		13'b1011100001001: color_data = 12'b001110100111;
		13'b1011100001010: color_data = 12'b001110100111;
		13'b1011100001011: color_data = 12'b001110100111;
		13'b1011100010011: color_data = 12'b001110100111;
		13'b1011100010100: color_data = 12'b001110100111;
		13'b1011100010101: color_data = 12'b001110100111;
		13'b1011100010110: color_data = 12'b001110100111;
		13'b1011100010111: color_data = 12'b001110100111;
		13'b1011100011000: color_data = 12'b001110100111;
		13'b1011100011001: color_data = 12'b001110100111;
		13'b1011100011010: color_data = 12'b001110100111;
		13'b1011100011011: color_data = 12'b001110100111;
		13'b1011100100000: color_data = 12'b001110100111;
		13'b1011100100001: color_data = 12'b001110100111;
		13'b1011100100010: color_data = 12'b001110100111;
		13'b1011100100011: color_data = 12'b001110100111;
		13'b1011100101011: color_data = 12'b001110100111;
		13'b1011100101100: color_data = 12'b001110100111;
		13'b1011100101101: color_data = 12'b001110100111;
		13'b1011100101110: color_data = 12'b001110100111;
		13'b1011100101111: color_data = 12'b001110100111;
		13'b1011100110000: color_data = 12'b001110100111;
		13'b1011100110101: color_data = 12'b001110100111;
		13'b1011100110110: color_data = 12'b001110100111;
		13'b1011100110111: color_data = 12'b001110100111;
		13'b1011100111000: color_data = 12'b001110100111;
		13'b1011100111001: color_data = 12'b001110100111;
		13'b1011100111010: color_data = 12'b001110100111;
		13'b1011100111011: color_data = 12'b001110100111;
		13'b1011100111100: color_data = 12'b001110100111;
		13'b1011100111101: color_data = 12'b001110100111;
		13'b1011100111110: color_data = 12'b001110100111;
		13'b1011101000011: color_data = 12'b001110100111;
		13'b1011101000100: color_data = 12'b001110100111;
		13'b1011101000101: color_data = 12'b001110100111;
		13'b1011101000110: color_data = 12'b001110100111;
		13'b1011101001000: color_data = 12'b001110100111;
		13'b1011101001001: color_data = 12'b001110100111;
		13'b1011101001010: color_data = 12'b001110100111;
		13'b1011101001011: color_data = 12'b001110100111;
		13'b1011101010011: color_data = 12'b001110100111;
		13'b1011101010100: color_data = 12'b001110100111;
		13'b1011101010101: color_data = 12'b001110100111;
		13'b1011101010110: color_data = 12'b001110100111;
		13'b1011101010111: color_data = 12'b001110100111;
		13'b1011101011000: color_data = 12'b001110100111;
		13'b1011101011101: color_data = 12'b001110100111;
		13'b1011101011110: color_data = 12'b001110100111;
		13'b1011101011111: color_data = 12'b001110100111;
		13'b1011101100000: color_data = 12'b001110100111;
		13'b1011101100001: color_data = 12'b001110100111;
		13'b1011101100010: color_data = 12'b001110100111;
		13'b1011101100011: color_data = 12'b001110100111;
		13'b1011101100100: color_data = 12'b001110100111;
		13'b1011101100101: color_data = 12'b001110100111;
		13'b1011101101010: color_data = 12'b001110100111;
		13'b1011101101011: color_data = 12'b001110100111;
		13'b1011101101100: color_data = 12'b001110100111;
		13'b1011101101101: color_data = 12'b001110100111;
		13'b1011101101110: color_data = 12'b001110100111;
		13'b1011101101111: color_data = 12'b001110100111;
		13'b1011101110000: color_data = 12'b001110100111;
		13'b1011101110001: color_data = 12'b001110100111;
		13'b1011101110010: color_data = 12'b001110100111;
		13'b1011101110011: color_data = 12'b001110100111;
		13'b1011101110100: color_data = 12'b001110100111;
		13'b1011101110101: color_data = 12'b001110100111;
		13'b1011101110110: color_data = 12'b001110100111;
		13'b1011101111111: color_data = 12'b001110100111;
		13'b1011110000000: color_data = 12'b001110100111;
		13'b1011110000001: color_data = 12'b001110100111;
		13'b1011110000010: color_data = 12'b001110100111;
		13'b1011110000011: color_data = 12'b001110100111;

		default: color_data = 12'b000000000000;
	endcase
endmodule
