`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.01.2025 14:38:02
// Design Name: 
// Module Name: lives_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lives_rom
	(
		input wire clk,
		input wire [3:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [3:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
	10'b0000000000: color_data = 12'b001110100111;
		10'b0000000001: color_data = 12'b001110100111;
		10'b0000000010: color_data = 12'b001110100111;
		10'b0000001100: color_data = 12'b001110100111;
		10'b0000001101: color_data = 12'b001110100111;
		10'b0000010001: color_data = 12'b001110100111;
		10'b0000010010: color_data = 12'b001110100111;
		10'b0000010111: color_data = 12'b001110100111;
		10'b0000011000: color_data = 12'b001110100111;
		10'b0000011001: color_data = 12'b001110100111;
		10'b0000011100: color_data = 12'b001110100111;
		10'b0000011101: color_data = 12'b001110100111;
		10'b0000011110: color_data = 12'b001110100111;
		10'b0000011111: color_data = 12'b001110100111;
		10'b0000100000: color_data = 12'b001110100111;
		10'b0000100001: color_data = 12'b001110100111;
		10'b0000100010: color_data = 12'b001110100111;
		10'b0000100011: color_data = 12'b001110100111;
		10'b0000100100: color_data = 12'b001110100111;
		10'b0000100111: color_data = 12'b001110100111;
		10'b0000101000: color_data = 12'b001110100111;
		10'b0000101001: color_data = 12'b001110100111;
		10'b0000101010: color_data = 12'b001110100111;
		10'b0000101011: color_data = 12'b001110100111;
		10'b0000101100: color_data = 12'b001110100111;
		10'b0000101101: color_data = 12'b001110100111;
		10'b0000101110: color_data = 12'b001110100111;
		10'b0000101111: color_data = 12'b001110100111;
		10'b0000110000: color_data = 12'b001110100111;
		10'b0001000000: color_data = 12'b001110100111;
		10'b0001000001: color_data = 12'b001110100111;
		10'b0001000010: color_data = 12'b001110100111;
		10'b0001001100: color_data = 12'b001110100111;
		10'b0001001101: color_data = 12'b001110100111;
		10'b0001010001: color_data = 12'b001110100111;
		10'b0001010010: color_data = 12'b001110100111;
		10'b0001010111: color_data = 12'b001110100111;
		10'b0001011000: color_data = 12'b001110100111;
		10'b0001011001: color_data = 12'b001110100111;
		10'b0001011100: color_data = 12'b001110100111;
		10'b0001011101: color_data = 12'b001110100111;
		10'b0001011110: color_data = 12'b001110100111;
		10'b0001011111: color_data = 12'b001110100111;
		10'b0001100000: color_data = 12'b001110100111;
		10'b0001100001: color_data = 12'b001110100111;
		10'b0001100010: color_data = 12'b001110100111;
		10'b0001100011: color_data = 12'b001110100111;
		10'b0001100100: color_data = 12'b001110100111;
		10'b0001100111: color_data = 12'b001110100111;
		10'b0001101000: color_data = 12'b001110100111;
		10'b0001101001: color_data = 12'b001110100111;
		10'b0001101010: color_data = 12'b001110100111;
		10'b0001101011: color_data = 12'b001110100111;
		10'b0001101100: color_data = 12'b001110100111;
		10'b0001101101: color_data = 12'b001110100111;
		10'b0001101110: color_data = 12'b001110100111;
		10'b0001101111: color_data = 12'b001110100111;
		10'b0001110000: color_data = 12'b001110100111;
		10'b0010000000: color_data = 12'b001110100111;
		10'b0010000001: color_data = 12'b001110100111;
		10'b0010000010: color_data = 12'b001110100111;
		10'b0010001100: color_data = 12'b001110100111;
		10'b0010001101: color_data = 12'b001110100111;
		10'b0010010001: color_data = 12'b001110100111;
		10'b0010010010: color_data = 12'b001110100111;
		10'b0010010111: color_data = 12'b001110100111;
		10'b0010011000: color_data = 12'b001110100111;
		10'b0010011001: color_data = 12'b001110100111;
		10'b0010011100: color_data = 12'b001110100111;
		10'b0010011101: color_data = 12'b001110100111;
		10'b0010011110: color_data = 12'b001110100111;
		10'b0010011111: color_data = 12'b001110100111;
		10'b0010100000: color_data = 12'b001110100111;
		10'b0010100001: color_data = 12'b001110100111;
		10'b0010100010: color_data = 12'b001110100111;
		10'b0010100011: color_data = 12'b001110100111;
		10'b0010100100: color_data = 12'b001110100111;
		10'b0010100111: color_data = 12'b001110100111;
		10'b0010101000: color_data = 12'b001110100111;
		10'b0010101001: color_data = 12'b001110100111;
		10'b0010101010: color_data = 12'b001110100111;
		10'b0010101011: color_data = 12'b001110100111;
		10'b0010101100: color_data = 12'b001110100111;
		10'b0010101101: color_data = 12'b001110100111;
		10'b0010101110: color_data = 12'b001110100111;
		10'b0010101111: color_data = 12'b001110100111;
		10'b0010110000: color_data = 12'b001110100111;
		10'b0010110101: color_data = 12'b001110100111;
		10'b0010110110: color_data = 12'b001110100111;
		10'b0010110111: color_data = 12'b001110100111;
		10'b0011000000: color_data = 12'b001110100111;
		10'b0011000001: color_data = 12'b001110100111;
		10'b0011000010: color_data = 12'b001110100111;
		10'b0011001100: color_data = 12'b001110100111;
		10'b0011001101: color_data = 12'b001110100111;
		10'b0011010001: color_data = 12'b001110100111;
		10'b0011010010: color_data = 12'b001110100111;
		10'b0011010111: color_data = 12'b001110100111;
		10'b0011011000: color_data = 12'b001110100111;
		10'b0011011001: color_data = 12'b001110100111;
		10'b0011011100: color_data = 12'b001110100111;
		10'b0011011101: color_data = 12'b001110100111;
		10'b0011100111: color_data = 12'b001110100111;
		10'b0011101000: color_data = 12'b001110100111;
		10'b0011101001: color_data = 12'b001110100111;
		10'b0011110101: color_data = 12'b001110100111;
		10'b0011110110: color_data = 12'b001110100111;
		10'b0011110111: color_data = 12'b001110100111;
		10'b0100000000: color_data = 12'b001110100111;
		10'b0100000001: color_data = 12'b001110100111;
		10'b0100000010: color_data = 12'b001110100111;
		10'b0100001100: color_data = 12'b001110100111;
		10'b0100001101: color_data = 12'b001110100111;
		10'b0100010001: color_data = 12'b001110100111;
		10'b0100010010: color_data = 12'b001110100111;
		10'b0100010111: color_data = 12'b001110100111;
		10'b0100011000: color_data = 12'b001110100111;
		10'b0100011001: color_data = 12'b001110100111;
		10'b0100011100: color_data = 12'b001110100111;
		10'b0100011101: color_data = 12'b001110100111;
		10'b0100100111: color_data = 12'b001110100111;
		10'b0100101000: color_data = 12'b001110100111;
		10'b0100101001: color_data = 12'b001110100111;
		10'b0100110101: color_data = 12'b001110100111;
		10'b0100110110: color_data = 12'b001110100111;
		10'b0100110111: color_data = 12'b001110100111;
		10'b0101000000: color_data = 12'b001110100111;
		10'b0101000001: color_data = 12'b001110100111;
		10'b0101000010: color_data = 12'b001110100111;
		10'b0101001100: color_data = 12'b001110100111;
		10'b0101001101: color_data = 12'b001110100111;
		10'b0101010001: color_data = 12'b001110100111;
		10'b0101010010: color_data = 12'b001110100111;
		10'b0101010111: color_data = 12'b001110100111;
		10'b0101011000: color_data = 12'b001110100111;
		10'b0101011001: color_data = 12'b001110100111;
		10'b0101011100: color_data = 12'b001110100111;
		10'b0101011101: color_data = 12'b001110100111;
		10'b0101011110: color_data = 12'b001110100111;
		10'b0101011111: color_data = 12'b001110100111;
		10'b0101100000: color_data = 12'b001110100111;
		10'b0101100001: color_data = 12'b001110100111;
		10'b0101100010: color_data = 12'b001110100111;
		10'b0101100011: color_data = 12'b001110100111;
		10'b0101100100: color_data = 12'b001110100111;
		10'b0101100111: color_data = 12'b001110100111;
		10'b0101101000: color_data = 12'b001110100111;
		10'b0101101001: color_data = 12'b001110100111;
		10'b0101101010: color_data = 12'b001110100111;
		10'b0101101011: color_data = 12'b001110100111;
		10'b0101101100: color_data = 12'b001110100111;
		10'b0101101101: color_data = 12'b001110100111;
		10'b0101101110: color_data = 12'b001110100111;
		10'b0101101111: color_data = 12'b001110100111;
		10'b0101110000: color_data = 12'b001110100111;
		10'b0110000000: color_data = 12'b001110100111;
		10'b0110000001: color_data = 12'b001110100111;
		10'b0110000010: color_data = 12'b001110100111;
		10'b0110001100: color_data = 12'b001110100111;
		10'b0110001101: color_data = 12'b001110100111;
		10'b0110010001: color_data = 12'b001110100111;
		10'b0110010010: color_data = 12'b001110100111;
		10'b0110010111: color_data = 12'b001110100111;
		10'b0110011000: color_data = 12'b001110100111;
		10'b0110011001: color_data = 12'b001110100111;
		10'b0110011100: color_data = 12'b001110100111;
		10'b0110011101: color_data = 12'b001110100111;
		10'b0110011110: color_data = 12'b001110100111;
		10'b0110011111: color_data = 12'b001110100111;
		10'b0110100000: color_data = 12'b001110100111;
		10'b0110100001: color_data = 12'b001110100111;
		10'b0110100010: color_data = 12'b001110100111;
		10'b0110100011: color_data = 12'b001110100111;
		10'b0110100100: color_data = 12'b001110100111;
		10'b0110100111: color_data = 12'b001110100111;
		10'b0110101000: color_data = 12'b001110100111;
		10'b0110101001: color_data = 12'b001110100111;
		10'b0110101010: color_data = 12'b001110100111;
		10'b0110101011: color_data = 12'b001110100111;
		10'b0110101100: color_data = 12'b001110100111;
		10'b0110101101: color_data = 12'b001110100111;
		10'b0110101110: color_data = 12'b001110100111;
		10'b0110101111: color_data = 12'b001110100111;
		10'b0110110000: color_data = 12'b001110100111;
		10'b0111000000: color_data = 12'b001110100111;
		10'b0111000001: color_data = 12'b001110100111;
		10'b0111000010: color_data = 12'b001110100111;
		10'b0111001100: color_data = 12'b001110100111;
		10'b0111001101: color_data = 12'b001110100111;
		10'b0111010001: color_data = 12'b001110100111;
		10'b0111010010: color_data = 12'b001110100111;
		10'b0111010111: color_data = 12'b001110100111;
		10'b0111011000: color_data = 12'b001110100111;
		10'b0111011001: color_data = 12'b001110100111;
		10'b0111011100: color_data = 12'b001110100111;
		10'b0111011101: color_data = 12'b001110100111;
		10'b0111011110: color_data = 12'b001110100111;
		10'b0111011111: color_data = 12'b001110100111;
		10'b0111100000: color_data = 12'b001110100111;
		10'b0111100001: color_data = 12'b001110100111;
		10'b0111100010: color_data = 12'b001110100111;
		10'b0111100011: color_data = 12'b001110100111;
		10'b0111100100: color_data = 12'b001110100111;
		10'b0111100111: color_data = 12'b001110100111;
		10'b0111101000: color_data = 12'b001110100111;
		10'b0111101001: color_data = 12'b001110100111;
		10'b0111101010: color_data = 12'b001110100111;
		10'b0111101011: color_data = 12'b001110100111;
		10'b0111101100: color_data = 12'b001110100111;
		10'b0111101101: color_data = 12'b001110100111;
		10'b0111101110: color_data = 12'b001110100111;
		10'b0111101111: color_data = 12'b001110100111;
		10'b0111110000: color_data = 12'b001110100111;
		10'b1000000000: color_data = 12'b001110100111;
		10'b1000000001: color_data = 12'b001110100111;
		10'b1000000010: color_data = 12'b001110100111;
		10'b1000001100: color_data = 12'b001110100111;
		10'b1000001101: color_data = 12'b001110100111;
		10'b1000010001: color_data = 12'b001110100111;
		10'b1000010010: color_data = 12'b001110100111;
		10'b1000010111: color_data = 12'b001110100111;
		10'b1000011000: color_data = 12'b001110100111;
		10'b1000011001: color_data = 12'b001110100111;
		10'b1000011100: color_data = 12'b001110100111;
		10'b1000011101: color_data = 12'b001110100111;
		10'b1000101110: color_data = 12'b001110100111;
		10'b1000101111: color_data = 12'b001110100111;
		10'b1000110000: color_data = 12'b001110100111;
		10'b1000110101: color_data = 12'b001110100111;
		10'b1000110110: color_data = 12'b001110100111;
		10'b1000110111: color_data = 12'b001110100111;
		10'b1001000000: color_data = 12'b001110100111;
		10'b1001000001: color_data = 12'b001110100111;
		10'b1001000010: color_data = 12'b001110100111;
		10'b1001001100: color_data = 12'b001110100111;
		10'b1001001101: color_data = 12'b001110100111;
		10'b1001010001: color_data = 12'b001110100111;
		10'b1001010010: color_data = 12'b001110100111;
		10'b1001010111: color_data = 12'b001110100111;
		10'b1001011000: color_data = 12'b001110100111;
		10'b1001011001: color_data = 12'b001110100111;
		10'b1001011100: color_data = 12'b001110100111;
		10'b1001011101: color_data = 12'b001110100111;
		10'b1001101110: color_data = 12'b001110100111;
		10'b1001101111: color_data = 12'b001110100111;
		10'b1001110000: color_data = 12'b001110100111;
		10'b1001110101: color_data = 12'b001110100111;
		10'b1001110110: color_data = 12'b001110100111;
		10'b1001110111: color_data = 12'b001110100111;
		10'b1010000000: color_data = 12'b001110100111;
		10'b1010000001: color_data = 12'b001110100111;
		10'b1010000010: color_data = 12'b001110100111;
		10'b1010001100: color_data = 12'b001110100111;
		10'b1010001101: color_data = 12'b001110100111;
		10'b1010010001: color_data = 12'b001110100111;
		10'b1010010010: color_data = 12'b001110100111;
		10'b1010010111: color_data = 12'b001110100111;
		10'b1010011000: color_data = 12'b001110100111;
		10'b1010011001: color_data = 12'b001110100111;
		10'b1010011100: color_data = 12'b001110100111;
		10'b1010011101: color_data = 12'b001110100111;
		10'b1010101110: color_data = 12'b001110100111;
		10'b1010101111: color_data = 12'b001110100111;
		10'b1010110000: color_data = 12'b001110100111;
		10'b1010110101: color_data = 12'b001110100111;
		10'b1010110110: color_data = 12'b001110100111;
		10'b1010110111: color_data = 12'b001110100111;
		10'b1011000000: color_data = 12'b001110100111;
		10'b1011000001: color_data = 12'b001110100111;
		10'b1011000010: color_data = 12'b001110100111;
		10'b1011000011: color_data = 12'b001110100111;
		10'b1011000100: color_data = 12'b001110100111;
		10'b1011000101: color_data = 12'b001110100111;
		10'b1011000110: color_data = 12'b001110100111;
		10'b1011000111: color_data = 12'b001110100111;
		10'b1011001000: color_data = 12'b001110100111;
		10'b1011001001: color_data = 12'b001110100111;
		10'b1011001100: color_data = 12'b001110100111;
		10'b1011001101: color_data = 12'b001110100111;
		10'b1011010001: color_data = 12'b001110100111;
		10'b1011010010: color_data = 12'b001110100111;
		10'b1011010011: color_data = 12'b001110100111;
		10'b1011010100: color_data = 12'b001110100111;
		10'b1011010101: color_data = 12'b001110100111;
		10'b1011010110: color_data = 12'b001110100111;
		10'b1011011100: color_data = 12'b001110100111;
		10'b1011011101: color_data = 12'b001110100111;
		10'b1011011110: color_data = 12'b001110100111;
		10'b1011011111: color_data = 12'b001110100111;
		10'b1011100000: color_data = 12'b001110100111;
		10'b1011100001: color_data = 12'b001110100111;
		10'b1011100010: color_data = 12'b001110100111;
		10'b1011100011: color_data = 12'b001110100111;
		10'b1011100100: color_data = 12'b001110100111;
		10'b1011100111: color_data = 12'b001110100111;
		10'b1011101000: color_data = 12'b001110100111;
		10'b1011101001: color_data = 12'b001110100111;
		10'b1011101010: color_data = 12'b001110100111;
		10'b1011101011: color_data = 12'b001110100111;
		10'b1011101100: color_data = 12'b001110100111;
		10'b1011101101: color_data = 12'b001110100111;
		10'b1011101110: color_data = 12'b001110100111;
		10'b1011101111: color_data = 12'b001110100111;
		10'b1011110000: color_data = 12'b001110100111;
		10'b1100000000: color_data = 12'b001110100111;
		10'b1100000001: color_data = 12'b001110100111;
		10'b1100000010: color_data = 12'b001110100111;
		10'b1100000011: color_data = 12'b001110100111;
		10'b1100000100: color_data = 12'b001110100111;
		10'b1100000101: color_data = 12'b001110100111;
		10'b1100000110: color_data = 12'b001110100111;
		10'b1100000111: color_data = 12'b001110100111;
		10'b1100001000: color_data = 12'b001110100111;
		10'b1100001001: color_data = 12'b001110100111;
		10'b1100001100: color_data = 12'b001110100111;
		10'b1100001101: color_data = 12'b001110100111;
		10'b1100010001: color_data = 12'b001110100111;
		10'b1100010010: color_data = 12'b001110100111;
		10'b1100010011: color_data = 12'b001110100111;
		10'b1100010100: color_data = 12'b001110100111;
		10'b1100010101: color_data = 12'b001110100111;
		10'b1100010110: color_data = 12'b001110100111;
		10'b1100011100: color_data = 12'b001110100111;
		10'b1100011101: color_data = 12'b001110100111;
		10'b1100011110: color_data = 12'b001110100111;
		10'b1100011111: color_data = 12'b001110100111;
		10'b1100100000: color_data = 12'b001110100111;
		10'b1100100001: color_data = 12'b001110100111;
		10'b1100100010: color_data = 12'b001110100111;
		10'b1100100011: color_data = 12'b001110100111;
		10'b1100100100: color_data = 12'b001110100111;
		10'b1100100111: color_data = 12'b001110100111;
		10'b1100101000: color_data = 12'b001110100111;
		10'b1100101001: color_data = 12'b001110100111;
		10'b1100101010: color_data = 12'b001110100111;
		10'b1100101011: color_data = 12'b001110100111;
		10'b1100101100: color_data = 12'b001110100111;
		10'b1100101101: color_data = 12'b001110100111;
		10'b1100101110: color_data = 12'b001110100111;
		10'b1100101111: color_data = 12'b001110100111;
		10'b1100110000: color_data = 12'b001110100111;

		default: color_data = 12'b000000000000;
	endcase
endmodule
