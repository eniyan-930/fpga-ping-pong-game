`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.01.2025 17:07:59
// Design Name: 
// Module Name: multi_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module multi_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
        14'b00000000000000: color_data = 12'b110011110111;
		14'b00000000000001: color_data = 12'b110011110111;
		14'b00000000000010: color_data = 12'b110011110111;
		14'b00000000000011: color_data = 12'b110011110111;
		14'b00000000000100: color_data = 12'b110011110111;
		14'b00000000000101: color_data = 12'b110011110111;
		14'b00000000000110: color_data = 12'b110011110111;
		14'b00000000000111: color_data = 12'b110011110111;
		14'b00000000001000: color_data = 12'b110011110111;
		14'b00000000001001: color_data = 12'b110011110111;
		14'b00000000001010: color_data = 12'b110011110111;
		14'b00000000001011: color_data = 12'b110011110111;
		14'b00000000001100: color_data = 12'b110011110111;
		14'b00000000001101: color_data = 12'b110011110111;
		14'b00000000001110: color_data = 12'b110011110111;
		14'b00000000001111: color_data = 12'b110011110111;
		14'b00000000010000: color_data = 12'b110011110111;
		14'b00000000010001: color_data = 12'b110011110111;
		14'b00000000010010: color_data = 12'b110011110111;
		14'b00000000010011: color_data = 12'b110011110111;
		14'b00000000010100: color_data = 12'b110011110111;
		14'b00000000010101: color_data = 12'b110011110111;
		14'b00000000010110: color_data = 12'b110011110111;
		14'b00000000010111: color_data = 12'b110011110111;
		14'b00000000011000: color_data = 12'b110011110111;
		14'b00000000011001: color_data = 12'b110011110111;
		14'b00000000011010: color_data = 12'b110011110111;
		14'b00000000110110: color_data = 12'b110011110111;
		14'b00000000110111: color_data = 12'b110011110111;
		14'b00000000111000: color_data = 12'b110011110111;
		14'b00000000111001: color_data = 12'b110011110111;
		14'b00000000111010: color_data = 12'b110011110111;
		14'b00000000111011: color_data = 12'b110011110111;
		14'b00000001000001: color_data = 12'b110011110111;
		14'b00000001000010: color_data = 12'b110011110111;
		14'b00000001000011: color_data = 12'b110011110111;
		14'b00000001000100: color_data = 12'b110011110111;
		14'b00000001000101: color_data = 12'b110011110111;
		14'b00000001010001: color_data = 12'b110011110111;
		14'b00000001010010: color_data = 12'b110011110111;
		14'b00000001010011: color_data = 12'b110011110111;
		14'b00000001010100: color_data = 12'b110011110111;
		14'b00000001010101: color_data = 12'b110011110111;
		14'b00000001010110: color_data = 12'b110011110111;
		14'b00000001100001: color_data = 12'b110011110111;
		14'b00000001100010: color_data = 12'b110011110111;
		14'b00000001100011: color_data = 12'b110011110111;
		14'b00000001100100: color_data = 12'b110011110111;
		14'b00000001100101: color_data = 12'b110011110111;
		14'b00000001100110: color_data = 12'b110011110111;
		14'b00000001100111: color_data = 12'b110011110111;
		14'b00000001101000: color_data = 12'b110011110111;
		14'b00000001101001: color_data = 12'b110011110111;
		14'b00000001101010: color_data = 12'b110011110111;
		14'b00000001101011: color_data = 12'b110011110111;
		14'b00000001101100: color_data = 12'b110011110111;
		14'b00000001101101: color_data = 12'b110011110111;
		14'b00000001101110: color_data = 12'b110011110111;
		14'b00000001101111: color_data = 12'b110011110111;
		14'b00000001110000: color_data = 12'b110011110111;
		14'b00000001110001: color_data = 12'b110011110111;
		14'b00000001110010: color_data = 12'b110011110111;
		14'b00000001110011: color_data = 12'b110011110111;
		14'b00000001110100: color_data = 12'b110011110111;
		14'b00000001110101: color_data = 12'b110011110111;
		14'b00000001110110: color_data = 12'b110011110111;
		14'b00000001111100: color_data = 12'b110011110111;
		14'b00000001111101: color_data = 12'b110011110111;
		14'b00000001111110: color_data = 12'b110011110111;
		14'b00000001111111: color_data = 12'b110011110111;
		14'b00000010000000: color_data = 12'b110011110111;
		14'b00000010000001: color_data = 12'b110011110111;
		14'b00000100000000: color_data = 12'b110011110111;
		14'b00000100000001: color_data = 12'b110011110111;
		14'b00000100000010: color_data = 12'b110011110111;
		14'b00000100000011: color_data = 12'b110011110111;
		14'b00000100000100: color_data = 12'b110011110111;
		14'b00000100000101: color_data = 12'b110011110111;
		14'b00000100000110: color_data = 12'b110011110111;
		14'b00000100000111: color_data = 12'b110011110111;
		14'b00000100001000: color_data = 12'b110011110111;
		14'b00000100001001: color_data = 12'b110011110111;
		14'b00000100001010: color_data = 12'b110011110111;
		14'b00000100001011: color_data = 12'b110011110111;
		14'b00000100001100: color_data = 12'b110011110111;
		14'b00000100001101: color_data = 12'b110011110111;
		14'b00000100001110: color_data = 12'b110011110111;
		14'b00000100001111: color_data = 12'b110011110111;
		14'b00000100010000: color_data = 12'b110011110111;
		14'b00000100010001: color_data = 12'b110011110111;
		14'b00000100010010: color_data = 12'b110011110111;
		14'b00000100010011: color_data = 12'b110011110111;
		14'b00000100010100: color_data = 12'b110011110111;
		14'b00000100010101: color_data = 12'b110011110111;
		14'b00000100010110: color_data = 12'b110011110111;
		14'b00000100010111: color_data = 12'b110011110111;
		14'b00000100011000: color_data = 12'b110011110111;
		14'b00000100011001: color_data = 12'b110011110111;
		14'b00000100011010: color_data = 12'b110011110111;
		14'b00000100110110: color_data = 12'b110011110111;
		14'b00000100110111: color_data = 12'b110011110111;
		14'b00000100111000: color_data = 12'b110011110111;
		14'b00000100111001: color_data = 12'b110011110111;
		14'b00000100111010: color_data = 12'b110011110111;
		14'b00000100111011: color_data = 12'b110011110111;
		14'b00000101000001: color_data = 12'b110011110111;
		14'b00000101000010: color_data = 12'b110011110111;
		14'b00000101000011: color_data = 12'b110011110111;
		14'b00000101000100: color_data = 12'b110011110111;
		14'b00000101000101: color_data = 12'b110011110111;
		14'b00000101010001: color_data = 12'b110011110111;
		14'b00000101010010: color_data = 12'b110011110111;
		14'b00000101010011: color_data = 12'b110011110111;
		14'b00000101010100: color_data = 12'b110011110111;
		14'b00000101010101: color_data = 12'b110011110111;
		14'b00000101010110: color_data = 12'b110011110111;
		14'b00000101100001: color_data = 12'b110011110111;
		14'b00000101100010: color_data = 12'b110011110111;
		14'b00000101100011: color_data = 12'b110011110111;
		14'b00000101100100: color_data = 12'b110011110111;
		14'b00000101100101: color_data = 12'b110011110111;
		14'b00000101100110: color_data = 12'b110011110111;
		14'b00000101100111: color_data = 12'b110011110111;
		14'b00000101101000: color_data = 12'b110011110111;
		14'b00000101101001: color_data = 12'b110011110111;
		14'b00000101101010: color_data = 12'b110011110111;
		14'b00000101101011: color_data = 12'b110011110111;
		14'b00000101101100: color_data = 12'b110011110111;
		14'b00000101101101: color_data = 12'b110011110111;
		14'b00000101101110: color_data = 12'b110011110111;
		14'b00000101101111: color_data = 12'b110011110111;
		14'b00000101110000: color_data = 12'b110011110111;
		14'b00000101110001: color_data = 12'b110011110111;
		14'b00000101110010: color_data = 12'b110011110111;
		14'b00000101110011: color_data = 12'b110011110111;
		14'b00000101110100: color_data = 12'b110011110111;
		14'b00000101110101: color_data = 12'b110011110111;
		14'b00000101110110: color_data = 12'b110011110111;
		14'b00000101111100: color_data = 12'b110011110111;
		14'b00000101111101: color_data = 12'b110011110111;
		14'b00000101111110: color_data = 12'b110011110111;
		14'b00000101111111: color_data = 12'b110011110111;
		14'b00000110000000: color_data = 12'b110011110111;
		14'b00000110000001: color_data = 12'b110011110111;
		14'b00001000000000: color_data = 12'b110011110111;
		14'b00001000000001: color_data = 12'b110011110111;
		14'b00001000000010: color_data = 12'b110011110111;
		14'b00001000000011: color_data = 12'b110011110111;
		14'b00001000000100: color_data = 12'b110011110111;
		14'b00001000000101: color_data = 12'b110011110111;
		14'b00001000000110: color_data = 12'b110011110111;
		14'b00001000000111: color_data = 12'b110011110111;
		14'b00001000001000: color_data = 12'b110011110111;
		14'b00001000001001: color_data = 12'b110011110111;
		14'b00001000001010: color_data = 12'b110011110111;
		14'b00001000001011: color_data = 12'b110011110111;
		14'b00001000001100: color_data = 12'b110011110111;
		14'b00001000001101: color_data = 12'b110011110111;
		14'b00001000001110: color_data = 12'b110011110111;
		14'b00001000001111: color_data = 12'b110011110111;
		14'b00001000010000: color_data = 12'b110011110111;
		14'b00001000010001: color_data = 12'b110011110111;
		14'b00001000010010: color_data = 12'b110011110111;
		14'b00001000010011: color_data = 12'b110011110111;
		14'b00001000010100: color_data = 12'b110011110111;
		14'b00001000010101: color_data = 12'b110011110111;
		14'b00001000010110: color_data = 12'b110011110111;
		14'b00001000010111: color_data = 12'b110011110111;
		14'b00001000011000: color_data = 12'b110011110111;
		14'b00001000011001: color_data = 12'b110011110111;
		14'b00001000011010: color_data = 12'b110011110111;
		14'b00001000110110: color_data = 12'b110011110111;
		14'b00001000110111: color_data = 12'b110011110111;
		14'b00001000111000: color_data = 12'b110011110111;
		14'b00001000111001: color_data = 12'b110011110111;
		14'b00001000111010: color_data = 12'b110011110111;
		14'b00001000111011: color_data = 12'b110011110111;
		14'b00001001000001: color_data = 12'b110011110111;
		14'b00001001000010: color_data = 12'b110011110111;
		14'b00001001000011: color_data = 12'b110011110111;
		14'b00001001000100: color_data = 12'b110011110111;
		14'b00001001000101: color_data = 12'b110011110111;
		14'b00001001010001: color_data = 12'b110011110111;
		14'b00001001010010: color_data = 12'b110011110111;
		14'b00001001010011: color_data = 12'b110011110111;
		14'b00001001010100: color_data = 12'b110011110111;
		14'b00001001010101: color_data = 12'b110011110111;
		14'b00001001010110: color_data = 12'b110011110111;
		14'b00001001100001: color_data = 12'b110011110111;
		14'b00001001100010: color_data = 12'b110011110111;
		14'b00001001100011: color_data = 12'b110011110111;
		14'b00001001100100: color_data = 12'b110011110111;
		14'b00001001100101: color_data = 12'b110011110111;
		14'b00001001100110: color_data = 12'b110011110111;
		14'b00001001100111: color_data = 12'b110011110111;
		14'b00001001101000: color_data = 12'b110011110111;
		14'b00001001101001: color_data = 12'b110011110111;
		14'b00001001101010: color_data = 12'b110011110111;
		14'b00001001101011: color_data = 12'b110011110111;
		14'b00001001101100: color_data = 12'b110011110111;
		14'b00001001101101: color_data = 12'b110011110111;
		14'b00001001101110: color_data = 12'b110011110111;
		14'b00001001101111: color_data = 12'b110011110111;
		14'b00001001110000: color_data = 12'b110011110111;
		14'b00001001110001: color_data = 12'b110011110111;
		14'b00001001110010: color_data = 12'b110011110111;
		14'b00001001110011: color_data = 12'b110011110111;
		14'b00001001110100: color_data = 12'b110011110111;
		14'b00001001110101: color_data = 12'b110011110111;
		14'b00001001110110: color_data = 12'b110011110111;
		14'b00001001111100: color_data = 12'b110011110111;
		14'b00001001111101: color_data = 12'b110011110111;
		14'b00001001111110: color_data = 12'b110011110111;
		14'b00001001111111: color_data = 12'b110011110111;
		14'b00001010000000: color_data = 12'b110011110111;
		14'b00001010000001: color_data = 12'b110011110111;
		14'b00001100000000: color_data = 12'b110011110111;
		14'b00001100000001: color_data = 12'b110011110111;
		14'b00001100000010: color_data = 12'b110011110111;
		14'b00001100000011: color_data = 12'b110011110111;
		14'b00001100000100: color_data = 12'b110011110111;
		14'b00001100000101: color_data = 12'b110011110111;
		14'b00001100000110: color_data = 12'b110011110111;
		14'b00001100000111: color_data = 12'b110011110111;
		14'b00001100001000: color_data = 12'b110011110111;
		14'b00001100001001: color_data = 12'b110011110111;
		14'b00001100001010: color_data = 12'b110011110111;
		14'b00001100001011: color_data = 12'b110011110111;
		14'b00001100001100: color_data = 12'b110011110111;
		14'b00001100001101: color_data = 12'b110011110111;
		14'b00001100001110: color_data = 12'b110011110111;
		14'b00001100001111: color_data = 12'b110011110111;
		14'b00001100010000: color_data = 12'b110011110111;
		14'b00001100010001: color_data = 12'b110011110111;
		14'b00001100010010: color_data = 12'b110011110111;
		14'b00001100010011: color_data = 12'b110011110111;
		14'b00001100010100: color_data = 12'b110011110111;
		14'b00001100010101: color_data = 12'b110011110111;
		14'b00001100010110: color_data = 12'b110011110111;
		14'b00001100010111: color_data = 12'b110011110111;
		14'b00001100011000: color_data = 12'b110011110111;
		14'b00001100011001: color_data = 12'b110011110111;
		14'b00001100011010: color_data = 12'b110011110111;
		14'b00001100110110: color_data = 12'b110011110111;
		14'b00001100110111: color_data = 12'b110011110111;
		14'b00001100111000: color_data = 12'b110011110111;
		14'b00001100111001: color_data = 12'b110011110111;
		14'b00001100111010: color_data = 12'b110011110111;
		14'b00001100111011: color_data = 12'b110011110111;
		14'b00001101000001: color_data = 12'b110011110111;
		14'b00001101000010: color_data = 12'b110011110111;
		14'b00001101000011: color_data = 12'b110011110111;
		14'b00001101000100: color_data = 12'b110011110111;
		14'b00001101000101: color_data = 12'b110011110111;
		14'b00001101010001: color_data = 12'b110011110111;
		14'b00001101010010: color_data = 12'b110011110111;
		14'b00001101010011: color_data = 12'b110011110111;
		14'b00001101010100: color_data = 12'b110011110111;
		14'b00001101010101: color_data = 12'b110011110111;
		14'b00001101010110: color_data = 12'b110011110111;
		14'b00001101100001: color_data = 12'b110011110111;
		14'b00001101100010: color_data = 12'b110011110111;
		14'b00001101100011: color_data = 12'b110011110111;
		14'b00001101100100: color_data = 12'b110011110111;
		14'b00001101100101: color_data = 12'b110011110111;
		14'b00001101100110: color_data = 12'b110011110111;
		14'b00001101100111: color_data = 12'b110011110111;
		14'b00001101101000: color_data = 12'b110011110111;
		14'b00001101101001: color_data = 12'b110011110111;
		14'b00001101101010: color_data = 12'b110011110111;
		14'b00001101101011: color_data = 12'b110011110111;
		14'b00001101101100: color_data = 12'b110011110111;
		14'b00001101101101: color_data = 12'b110011110111;
		14'b00001101101110: color_data = 12'b110011110111;
		14'b00001101101111: color_data = 12'b110011110111;
		14'b00001101110000: color_data = 12'b110011110111;
		14'b00001101110001: color_data = 12'b110011110111;
		14'b00001101110010: color_data = 12'b110011110111;
		14'b00001101110011: color_data = 12'b110011110111;
		14'b00001101110100: color_data = 12'b110011110111;
		14'b00001101110101: color_data = 12'b110011110111;
		14'b00001101110110: color_data = 12'b110011110111;
		14'b00001101111100: color_data = 12'b110011110111;
		14'b00001101111101: color_data = 12'b110011110111;
		14'b00001101111110: color_data = 12'b110011110111;
		14'b00001101111111: color_data = 12'b110011110111;
		14'b00001110000000: color_data = 12'b110011110111;
		14'b00001110000001: color_data = 12'b110011110111;
		14'b00010000000000: color_data = 12'b110011110111;
		14'b00010000000001: color_data = 12'b110011110111;
		14'b00010000000010: color_data = 12'b110011110111;
		14'b00010000000011: color_data = 12'b110011110111;
		14'b00010000000100: color_data = 12'b110011110111;
		14'b00010000000101: color_data = 12'b110011110111;
		14'b00010000000110: color_data = 12'b110011110111;
		14'b00010000000111: color_data = 12'b110011110111;
		14'b00010000001000: color_data = 12'b110011110111;
		14'b00010000001001: color_data = 12'b110011110111;
		14'b00010000001010: color_data = 12'b110011110111;
		14'b00010000001011: color_data = 12'b110011110111;
		14'b00010000001100: color_data = 12'b110011110111;
		14'b00010000001101: color_data = 12'b110011110111;
		14'b00010000001110: color_data = 12'b110011110111;
		14'b00010000001111: color_data = 12'b110011110111;
		14'b00010000010000: color_data = 12'b110011110111;
		14'b00010000010001: color_data = 12'b110011110111;
		14'b00010000010010: color_data = 12'b110011110111;
		14'b00010000010011: color_data = 12'b110011110111;
		14'b00010000010100: color_data = 12'b110011110111;
		14'b00010000010101: color_data = 12'b110011110111;
		14'b00010000010110: color_data = 12'b110011110111;
		14'b00010000010111: color_data = 12'b110011110111;
		14'b00010000011000: color_data = 12'b110011110111;
		14'b00010000011001: color_data = 12'b110011110111;
		14'b00010000011010: color_data = 12'b110011110111;
		14'b00010000110110: color_data = 12'b110011110111;
		14'b00010000110111: color_data = 12'b110011110111;
		14'b00010000111000: color_data = 12'b110011110111;
		14'b00010000111001: color_data = 12'b110011110111;
		14'b00010000111010: color_data = 12'b110011110111;
		14'b00010000111011: color_data = 12'b110011110111;
		14'b00010001000001: color_data = 12'b110011110111;
		14'b00010001000010: color_data = 12'b110011110111;
		14'b00010001000011: color_data = 12'b110011110111;
		14'b00010001000100: color_data = 12'b110011110111;
		14'b00010001000101: color_data = 12'b110011110111;
		14'b00010001010001: color_data = 12'b110011110111;
		14'b00010001010010: color_data = 12'b110011110111;
		14'b00010001010011: color_data = 12'b110011110111;
		14'b00010001010100: color_data = 12'b110011110111;
		14'b00010001010101: color_data = 12'b110011110111;
		14'b00010001010110: color_data = 12'b110011110111;
		14'b00010001100001: color_data = 12'b110011110111;
		14'b00010001100010: color_data = 12'b110011110111;
		14'b00010001100011: color_data = 12'b110011110111;
		14'b00010001100100: color_data = 12'b110011110111;
		14'b00010001100101: color_data = 12'b110011110111;
		14'b00010001100110: color_data = 12'b110011110111;
		14'b00010001100111: color_data = 12'b110011110111;
		14'b00010001101000: color_data = 12'b110011110111;
		14'b00010001101001: color_data = 12'b110011110111;
		14'b00010001101010: color_data = 12'b110011110111;
		14'b00010001101011: color_data = 12'b110011110111;
		14'b00010001101100: color_data = 12'b110011110111;
		14'b00010001101101: color_data = 12'b110011110111;
		14'b00010001101110: color_data = 12'b110011110111;
		14'b00010001101111: color_data = 12'b110011110111;
		14'b00010001110000: color_data = 12'b110011110111;
		14'b00010001110001: color_data = 12'b110011110111;
		14'b00010001110010: color_data = 12'b110011110111;
		14'b00010001110011: color_data = 12'b110011110111;
		14'b00010001110100: color_data = 12'b110011110111;
		14'b00010001110101: color_data = 12'b110011110111;
		14'b00010001110110: color_data = 12'b110011110111;
		14'b00010001111100: color_data = 12'b110011110111;
		14'b00010001111101: color_data = 12'b110011110111;
		14'b00010001111110: color_data = 12'b110011110111;
		14'b00010001111111: color_data = 12'b110011110111;
		14'b00010010000000: color_data = 12'b110011110111;
		14'b00010010000001: color_data = 12'b110011110111;
		14'b00010100000000: color_data = 12'b110011110111;
		14'b00010100000001: color_data = 12'b110011110111;
		14'b00010100000010: color_data = 12'b110011110111;
		14'b00010100000011: color_data = 12'b110011110111;
		14'b00010100000100: color_data = 12'b110011110111;
		14'b00010100000101: color_data = 12'b110011110111;
		14'b00010100001011: color_data = 12'b110011110111;
		14'b00010100001100: color_data = 12'b110011110111;
		14'b00010100001101: color_data = 12'b110011110111;
		14'b00010100001110: color_data = 12'b110011110111;
		14'b00010100001111: color_data = 12'b110011110111;
		14'b00010100010000: color_data = 12'b110011110111;
		14'b00010100010110: color_data = 12'b110011110111;
		14'b00010100010111: color_data = 12'b110011110111;
		14'b00010100011000: color_data = 12'b110011110111;
		14'b00010100011001: color_data = 12'b110011110111;
		14'b00010100011010: color_data = 12'b110011110111;
		14'b00010100110110: color_data = 12'b110011110111;
		14'b00010100110111: color_data = 12'b110011110111;
		14'b00010100111000: color_data = 12'b110011110111;
		14'b00010100111001: color_data = 12'b110011110111;
		14'b00010100111010: color_data = 12'b110011110111;
		14'b00010100111011: color_data = 12'b110011110111;
		14'b00010101000001: color_data = 12'b110011110111;
		14'b00010101000010: color_data = 12'b110011110111;
		14'b00010101000011: color_data = 12'b110011110111;
		14'b00010101000100: color_data = 12'b110011110111;
		14'b00010101000101: color_data = 12'b110011110111;
		14'b00010101100001: color_data = 12'b110011110111;
		14'b00010101100010: color_data = 12'b110011110111;
		14'b00010101100011: color_data = 12'b110011110111;
		14'b00010101100100: color_data = 12'b110011110111;
		14'b00010101100101: color_data = 12'b110011110111;
		14'b00010101100110: color_data = 12'b110011110111;
		14'b00010101110010: color_data = 12'b110011110111;
		14'b00010101110011: color_data = 12'b110011110111;
		14'b00010101110100: color_data = 12'b110011110111;
		14'b00010101110101: color_data = 12'b110011110111;
		14'b00010101110110: color_data = 12'b110011110111;
		14'b00010101111100: color_data = 12'b110011110111;
		14'b00010101111101: color_data = 12'b110011110111;
		14'b00010101111110: color_data = 12'b110011110111;
		14'b00010101111111: color_data = 12'b110011110111;
		14'b00010110000000: color_data = 12'b110011110111;
		14'b00010110000001: color_data = 12'b110011110111;
		14'b00011000000000: color_data = 12'b110011110111;
		14'b00011000000001: color_data = 12'b110011110111;
		14'b00011000000010: color_data = 12'b110011110111;
		14'b00011000000011: color_data = 12'b110011110111;
		14'b00011000000100: color_data = 12'b110011110111;
		14'b00011000000101: color_data = 12'b110011110111;
		14'b00011000001011: color_data = 12'b110011110111;
		14'b00011000001100: color_data = 12'b110011110111;
		14'b00011000001101: color_data = 12'b110011110111;
		14'b00011000001110: color_data = 12'b110011110111;
		14'b00011000001111: color_data = 12'b110011110111;
		14'b00011000010000: color_data = 12'b110011110111;
		14'b00011000010110: color_data = 12'b110011110111;
		14'b00011000010111: color_data = 12'b110011110111;
		14'b00011000011000: color_data = 12'b110011110111;
		14'b00011000011001: color_data = 12'b110011110111;
		14'b00011000011010: color_data = 12'b110011110111;
		14'b00011000110110: color_data = 12'b110011110111;
		14'b00011000110111: color_data = 12'b110011110111;
		14'b00011000111000: color_data = 12'b110011110111;
		14'b00011000111001: color_data = 12'b110011110111;
		14'b00011000111010: color_data = 12'b110011110111;
		14'b00011000111011: color_data = 12'b110011110111;
		14'b00011001000001: color_data = 12'b110011110111;
		14'b00011001000010: color_data = 12'b110011110111;
		14'b00011001000011: color_data = 12'b110011110111;
		14'b00011001000100: color_data = 12'b110011110111;
		14'b00011001000101: color_data = 12'b110011110111;
		14'b00011001100001: color_data = 12'b110011110111;
		14'b00011001100010: color_data = 12'b110011110111;
		14'b00011001100011: color_data = 12'b110011110111;
		14'b00011001100100: color_data = 12'b110011110111;
		14'b00011001100101: color_data = 12'b110011110111;
		14'b00011001100110: color_data = 12'b110011110111;
		14'b00011001110010: color_data = 12'b110011110111;
		14'b00011001110011: color_data = 12'b110011110111;
		14'b00011001110100: color_data = 12'b110011110111;
		14'b00011001110101: color_data = 12'b110011110111;
		14'b00011001110110: color_data = 12'b110011110111;
		14'b00011001111100: color_data = 12'b110011110111;
		14'b00011001111101: color_data = 12'b110011110111;
		14'b00011001111110: color_data = 12'b110011110111;
		14'b00011001111111: color_data = 12'b110011110111;
		14'b00011010000000: color_data = 12'b110011110111;
		14'b00011010000001: color_data = 12'b110011110111;
		14'b00011100000000: color_data = 12'b110011110111;
		14'b00011100000001: color_data = 12'b110011110111;
		14'b00011100000010: color_data = 12'b110011110111;
		14'b00011100000011: color_data = 12'b110011110111;
		14'b00011100000100: color_data = 12'b110011110111;
		14'b00011100000101: color_data = 12'b110011110111;
		14'b00011100001011: color_data = 12'b110011110111;
		14'b00011100001100: color_data = 12'b110011110111;
		14'b00011100001101: color_data = 12'b110011110111;
		14'b00011100001110: color_data = 12'b110011110111;
		14'b00011100001111: color_data = 12'b110011110111;
		14'b00011100010000: color_data = 12'b110011110111;
		14'b00011100010110: color_data = 12'b110011110111;
		14'b00011100010111: color_data = 12'b110011110111;
		14'b00011100011000: color_data = 12'b110011110111;
		14'b00011100011001: color_data = 12'b110011110111;
		14'b00011100011010: color_data = 12'b110011110111;
		14'b00011100110110: color_data = 12'b110011110111;
		14'b00011100110111: color_data = 12'b110011110111;
		14'b00011100111000: color_data = 12'b110011110111;
		14'b00011100111001: color_data = 12'b110011110111;
		14'b00011100111010: color_data = 12'b110011110111;
		14'b00011100111011: color_data = 12'b110011110111;
		14'b00011101000001: color_data = 12'b110011110111;
		14'b00011101000010: color_data = 12'b110011110111;
		14'b00011101000011: color_data = 12'b110011110111;
		14'b00011101000100: color_data = 12'b110011110111;
		14'b00011101000101: color_data = 12'b110011110111;
		14'b00011101100001: color_data = 12'b110011110111;
		14'b00011101100010: color_data = 12'b110011110111;
		14'b00011101100011: color_data = 12'b110011110111;
		14'b00011101100100: color_data = 12'b110011110111;
		14'b00011101100101: color_data = 12'b110011110111;
		14'b00011101100110: color_data = 12'b110011110111;
		14'b00011101110010: color_data = 12'b110011110111;
		14'b00011101110011: color_data = 12'b110011110111;
		14'b00011101110100: color_data = 12'b110011110111;
		14'b00011101110101: color_data = 12'b110011110111;
		14'b00011101110110: color_data = 12'b110011110111;
		14'b00011101111100: color_data = 12'b110011110111;
		14'b00011101111101: color_data = 12'b110011110111;
		14'b00011101111110: color_data = 12'b110011110111;
		14'b00011101111111: color_data = 12'b110011110111;
		14'b00011110000000: color_data = 12'b110011110111;
		14'b00011110000001: color_data = 12'b110011110111;
		14'b00100000000000: color_data = 12'b110011110111;
		14'b00100000000001: color_data = 12'b110011110111;
		14'b00100000000010: color_data = 12'b110011110111;
		14'b00100000000011: color_data = 12'b110011110111;
		14'b00100000000100: color_data = 12'b110011110111;
		14'b00100000000101: color_data = 12'b110011110111;
		14'b00100000001011: color_data = 12'b110011110111;
		14'b00100000001100: color_data = 12'b110011110111;
		14'b00100000001101: color_data = 12'b110011110111;
		14'b00100000001110: color_data = 12'b110011110111;
		14'b00100000001111: color_data = 12'b110011110111;
		14'b00100000010000: color_data = 12'b110011110111;
		14'b00100000010110: color_data = 12'b110011110111;
		14'b00100000010111: color_data = 12'b110011110111;
		14'b00100000011000: color_data = 12'b110011110111;
		14'b00100000011001: color_data = 12'b110011110111;
		14'b00100000011010: color_data = 12'b110011110111;
		14'b00100000110110: color_data = 12'b110011110111;
		14'b00100000110111: color_data = 12'b110011110111;
		14'b00100000111000: color_data = 12'b110011110111;
		14'b00100000111001: color_data = 12'b110011110111;
		14'b00100000111010: color_data = 12'b110011110111;
		14'b00100000111011: color_data = 12'b110011110111;
		14'b00100001000001: color_data = 12'b110011110111;
		14'b00100001000010: color_data = 12'b110011110111;
		14'b00100001000011: color_data = 12'b110011110111;
		14'b00100001000100: color_data = 12'b110011110111;
		14'b00100001000101: color_data = 12'b110011110111;
		14'b00100001100001: color_data = 12'b110011110111;
		14'b00100001100010: color_data = 12'b110011110111;
		14'b00100001100011: color_data = 12'b110011110111;
		14'b00100001100100: color_data = 12'b110011110111;
		14'b00100001100101: color_data = 12'b110011110111;
		14'b00100001100110: color_data = 12'b110011110111;
		14'b00100001110010: color_data = 12'b110011110111;
		14'b00100001110011: color_data = 12'b110011110111;
		14'b00100001110100: color_data = 12'b110011110111;
		14'b00100001110101: color_data = 12'b110011110111;
		14'b00100001110110: color_data = 12'b110011110111;
		14'b00100001111100: color_data = 12'b110011110111;
		14'b00100001111101: color_data = 12'b110011110111;
		14'b00100001111110: color_data = 12'b110011110111;
		14'b00100001111111: color_data = 12'b110011110111;
		14'b00100010000000: color_data = 12'b110011110111;
		14'b00100010000001: color_data = 12'b110011110111;
		14'b00100100000000: color_data = 12'b110011110111;
		14'b00100100000001: color_data = 12'b110011110111;
		14'b00100100000010: color_data = 12'b110011110111;
		14'b00100100000011: color_data = 12'b110011110111;
		14'b00100100000100: color_data = 12'b110011110111;
		14'b00100100000101: color_data = 12'b110011110111;
		14'b00100100001011: color_data = 12'b110011110111;
		14'b00100100001100: color_data = 12'b110011110111;
		14'b00100100001101: color_data = 12'b110011110111;
		14'b00100100001110: color_data = 12'b110011110111;
		14'b00100100001111: color_data = 12'b110011110111;
		14'b00100100010000: color_data = 12'b110011110111;
		14'b00100100010110: color_data = 12'b110011110111;
		14'b00100100010111: color_data = 12'b110011110111;
		14'b00100100011000: color_data = 12'b110011110111;
		14'b00100100011001: color_data = 12'b110011110111;
		14'b00100100011010: color_data = 12'b110011110111;
		14'b00100100100001: color_data = 12'b110011110111;
		14'b00100100100010: color_data = 12'b110011110111;
		14'b00100100100011: color_data = 12'b110011110111;
		14'b00100100100100: color_data = 12'b110011110111;
		14'b00100100100101: color_data = 12'b110011110111;
		14'b00100100101100: color_data = 12'b110011110111;
		14'b00100100101101: color_data = 12'b110011110111;
		14'b00100100101110: color_data = 12'b110011110111;
		14'b00100100101111: color_data = 12'b110011110111;
		14'b00100100110000: color_data = 12'b110011110111;
		14'b00100100110110: color_data = 12'b110011110111;
		14'b00100100110111: color_data = 12'b110011110111;
		14'b00100100111000: color_data = 12'b110011110111;
		14'b00100100111001: color_data = 12'b110011110111;
		14'b00100100111010: color_data = 12'b110011110111;
		14'b00100100111011: color_data = 12'b110011110111;
		14'b00100101000001: color_data = 12'b110011110111;
		14'b00100101000010: color_data = 12'b110011110111;
		14'b00100101000011: color_data = 12'b110011110111;
		14'b00100101000100: color_data = 12'b110011110111;
		14'b00100101000101: color_data = 12'b110011110111;
		14'b00100101000110: color_data = 12'b110011110111;
		14'b00100101000111: color_data = 12'b110011110111;
		14'b00100101001000: color_data = 12'b110011110111;
		14'b00100101001001: color_data = 12'b110011110111;
		14'b00100101001010: color_data = 12'b110011110111;
		14'b00100101001011: color_data = 12'b110011110111;
		14'b00100101010001: color_data = 12'b110011110111;
		14'b00100101010010: color_data = 12'b110011110111;
		14'b00100101010011: color_data = 12'b110011110111;
		14'b00100101010100: color_data = 12'b110011110111;
		14'b00100101010101: color_data = 12'b110011110111;
		14'b00100101010110: color_data = 12'b110011110111;
		14'b00100101100001: color_data = 12'b110011110111;
		14'b00100101100010: color_data = 12'b110011110111;
		14'b00100101100011: color_data = 12'b110011110111;
		14'b00100101100100: color_data = 12'b110011110111;
		14'b00100101100101: color_data = 12'b110011110111;
		14'b00100101100110: color_data = 12'b110011110111;
		14'b00100101100111: color_data = 12'b110011110111;
		14'b00100101101000: color_data = 12'b110011110111;
		14'b00100101101001: color_data = 12'b110011110111;
		14'b00100101101010: color_data = 12'b110011110111;
		14'b00100101101011: color_data = 12'b110011110111;
		14'b00100101101100: color_data = 12'b110011110111;
		14'b00100101101101: color_data = 12'b110011110111;
		14'b00100101101110: color_data = 12'b110011110111;
		14'b00100101101111: color_data = 12'b110011110111;
		14'b00100101110000: color_data = 12'b110011110111;
		14'b00100101110001: color_data = 12'b110011110111;
		14'b00100101110010: color_data = 12'b110011110111;
		14'b00100101110011: color_data = 12'b110011110111;
		14'b00100101110100: color_data = 12'b110011110111;
		14'b00100101110101: color_data = 12'b110011110111;
		14'b00100101110110: color_data = 12'b110011110111;
		14'b00100101111100: color_data = 12'b110011110111;
		14'b00100101111101: color_data = 12'b110011110111;
		14'b00100101111110: color_data = 12'b110011110111;
		14'b00100101111111: color_data = 12'b110011110111;
		14'b00100110000000: color_data = 12'b110011110111;
		14'b00100110000001: color_data = 12'b110011110111;
		14'b00100110001100: color_data = 12'b110011110111;
		14'b00100110001101: color_data = 12'b110011110111;
		14'b00100110001110: color_data = 12'b110011110111;
		14'b00100110001111: color_data = 12'b110011110111;
		14'b00100110010000: color_data = 12'b110011110111;
		14'b00100110010001: color_data = 12'b110011110111;
		14'b00100110010010: color_data = 12'b110011110111;
		14'b00100110010011: color_data = 12'b110011110111;
		14'b00100110010100: color_data = 12'b110011110111;
		14'b00100110010101: color_data = 12'b110011110111;
		14'b00100110010110: color_data = 12'b110011110111;
		14'b00100110011101: color_data = 12'b110011110111;
		14'b00100110011110: color_data = 12'b110011110111;
		14'b00100110011111: color_data = 12'b110011110111;
		14'b00100110100000: color_data = 12'b110011110111;
		14'b00100110100001: color_data = 12'b110011110111;
		14'b00100110100111: color_data = 12'b110011110111;
		14'b00100110101000: color_data = 12'b110011110111;
		14'b00100110101001: color_data = 12'b110011110111;
		14'b00100110101010: color_data = 12'b110011110111;
		14'b00100110101011: color_data = 12'b110011110111;
		14'b00100110101100: color_data = 12'b110011110111;
		14'b00100110110010: color_data = 12'b110011110111;
		14'b00100110110011: color_data = 12'b110011110111;
		14'b00100110110100: color_data = 12'b110011110111;
		14'b00100110110101: color_data = 12'b110011110111;
		14'b00100110110110: color_data = 12'b110011110111;
		14'b00100110110111: color_data = 12'b110011110111;
		14'b00100110111000: color_data = 12'b110011110111;
		14'b00100110111001: color_data = 12'b110011110111;
		14'b00100110111010: color_data = 12'b110011110111;
		14'b00100110111011: color_data = 12'b110011110111;
		14'b00100110111100: color_data = 12'b110011110111;
		14'b00100110111101: color_data = 12'b110011110111;
		14'b00100110111110: color_data = 12'b110011110111;
		14'b00100110111111: color_data = 12'b110011110111;
		14'b00100111000000: color_data = 12'b110011110111;
		14'b00100111000001: color_data = 12'b110011110111;
		14'b00100111001000: color_data = 12'b110011110111;
		14'b00100111001001: color_data = 12'b110011110111;
		14'b00100111001010: color_data = 12'b110011110111;
		14'b00100111001011: color_data = 12'b110011110111;
		14'b00100111001100: color_data = 12'b110011110111;
		14'b00100111001101: color_data = 12'b110011110111;
		14'b00100111001110: color_data = 12'b110011110111;
		14'b00100111001111: color_data = 12'b110011110111;
		14'b00100111010000: color_data = 12'b110011110111;
		14'b00100111010001: color_data = 12'b110011110111;
		14'b00101000000000: color_data = 12'b110011110111;
		14'b00101000000001: color_data = 12'b110011110111;
		14'b00101000000010: color_data = 12'b110011110111;
		14'b00101000000011: color_data = 12'b110011110111;
		14'b00101000000100: color_data = 12'b110011110111;
		14'b00101000000101: color_data = 12'b110011110111;
		14'b00101000001011: color_data = 12'b110011110111;
		14'b00101000001100: color_data = 12'b110011110111;
		14'b00101000001101: color_data = 12'b110011110111;
		14'b00101000001110: color_data = 12'b110011110111;
		14'b00101000001111: color_data = 12'b110011110111;
		14'b00101000010000: color_data = 12'b110011110111;
		14'b00101000010110: color_data = 12'b110011110111;
		14'b00101000010111: color_data = 12'b110011110111;
		14'b00101000011000: color_data = 12'b110011110111;
		14'b00101000011001: color_data = 12'b110011110111;
		14'b00101000011010: color_data = 12'b110011110111;
		14'b00101000100001: color_data = 12'b110011110111;
		14'b00101000100010: color_data = 12'b110011110111;
		14'b00101000100011: color_data = 12'b110011110111;
		14'b00101000100100: color_data = 12'b110011110111;
		14'b00101000100101: color_data = 12'b110011110111;
		14'b00101000101100: color_data = 12'b110011110111;
		14'b00101000101101: color_data = 12'b110011110111;
		14'b00101000101110: color_data = 12'b110011110111;
		14'b00101000101111: color_data = 12'b110011110111;
		14'b00101000110000: color_data = 12'b110011110111;
		14'b00101000110110: color_data = 12'b110011110111;
		14'b00101000110111: color_data = 12'b110011110111;
		14'b00101000111000: color_data = 12'b110011110111;
		14'b00101000111001: color_data = 12'b110011110111;
		14'b00101000111010: color_data = 12'b110011110111;
		14'b00101000111011: color_data = 12'b110011110111;
		14'b00101001000001: color_data = 12'b110011110111;
		14'b00101001000010: color_data = 12'b110011110111;
		14'b00101001000011: color_data = 12'b110011110111;
		14'b00101001000100: color_data = 12'b110011110111;
		14'b00101001000101: color_data = 12'b110011110111;
		14'b00101001000110: color_data = 12'b110011110111;
		14'b00101001000111: color_data = 12'b110011110111;
		14'b00101001001000: color_data = 12'b110011110111;
		14'b00101001001001: color_data = 12'b110011110111;
		14'b00101001001010: color_data = 12'b110011110111;
		14'b00101001001011: color_data = 12'b110011110111;
		14'b00101001010001: color_data = 12'b110011110111;
		14'b00101001010010: color_data = 12'b110011110111;
		14'b00101001010011: color_data = 12'b110011110111;
		14'b00101001010100: color_data = 12'b110011110111;
		14'b00101001010101: color_data = 12'b110011110111;
		14'b00101001010110: color_data = 12'b110011110111;
		14'b00101001100001: color_data = 12'b110011110111;
		14'b00101001100010: color_data = 12'b110011110111;
		14'b00101001100011: color_data = 12'b110011110111;
		14'b00101001100100: color_data = 12'b110011110111;
		14'b00101001100101: color_data = 12'b110011110111;
		14'b00101001100110: color_data = 12'b110011110111;
		14'b00101001100111: color_data = 12'b110011110111;
		14'b00101001101000: color_data = 12'b110011110111;
		14'b00101001101001: color_data = 12'b110011110111;
		14'b00101001101010: color_data = 12'b110011110111;
		14'b00101001101011: color_data = 12'b110011110111;
		14'b00101001101100: color_data = 12'b110011110111;
		14'b00101001101101: color_data = 12'b110011110111;
		14'b00101001101110: color_data = 12'b110011110111;
		14'b00101001101111: color_data = 12'b110011110111;
		14'b00101001110000: color_data = 12'b110011110111;
		14'b00101001110001: color_data = 12'b110011110111;
		14'b00101001110010: color_data = 12'b110011110111;
		14'b00101001110011: color_data = 12'b110011110111;
		14'b00101001110100: color_data = 12'b110011110111;
		14'b00101001110101: color_data = 12'b110011110111;
		14'b00101001110110: color_data = 12'b110011110111;
		14'b00101001111100: color_data = 12'b110011110111;
		14'b00101001111101: color_data = 12'b110011110111;
		14'b00101001111110: color_data = 12'b110011110111;
		14'b00101001111111: color_data = 12'b110011110111;
		14'b00101010000000: color_data = 12'b110011110111;
		14'b00101010000001: color_data = 12'b110011110111;
		14'b00101010001100: color_data = 12'b110011110111;
		14'b00101010001101: color_data = 12'b110011110111;
		14'b00101010001110: color_data = 12'b110011110111;
		14'b00101010001111: color_data = 12'b110011110111;
		14'b00101010010000: color_data = 12'b110011110111;
		14'b00101010010001: color_data = 12'b110011110111;
		14'b00101010010010: color_data = 12'b110011110111;
		14'b00101010010011: color_data = 12'b110011110111;
		14'b00101010010100: color_data = 12'b110011110111;
		14'b00101010010101: color_data = 12'b110011110111;
		14'b00101010010110: color_data = 12'b110011110111;
		14'b00101010011101: color_data = 12'b110011110111;
		14'b00101010011110: color_data = 12'b110011110111;
		14'b00101010011111: color_data = 12'b110011110111;
		14'b00101010100000: color_data = 12'b110011110111;
		14'b00101010100001: color_data = 12'b110011110111;
		14'b00101010100111: color_data = 12'b110011110111;
		14'b00101010101000: color_data = 12'b110011110111;
		14'b00101010101001: color_data = 12'b110011110111;
		14'b00101010101010: color_data = 12'b110011110111;
		14'b00101010101011: color_data = 12'b110011110111;
		14'b00101010101100: color_data = 12'b110011110111;
		14'b00101010110010: color_data = 12'b110011110111;
		14'b00101010110011: color_data = 12'b110011110111;
		14'b00101010110100: color_data = 12'b110011110111;
		14'b00101010110101: color_data = 12'b110011110111;
		14'b00101010110110: color_data = 12'b110011110111;
		14'b00101010110111: color_data = 12'b110011110111;
		14'b00101010111000: color_data = 12'b110011110111;
		14'b00101010111001: color_data = 12'b110011110111;
		14'b00101010111010: color_data = 12'b110011110111;
		14'b00101010111011: color_data = 12'b110011110111;
		14'b00101010111100: color_data = 12'b110011110111;
		14'b00101010111101: color_data = 12'b110011110111;
		14'b00101010111110: color_data = 12'b110011110111;
		14'b00101010111111: color_data = 12'b110011110111;
		14'b00101011000000: color_data = 12'b110011110111;
		14'b00101011000001: color_data = 12'b110011110111;
		14'b00101011001000: color_data = 12'b110011110111;
		14'b00101011001001: color_data = 12'b110011110111;
		14'b00101011001010: color_data = 12'b110011110111;
		14'b00101011001011: color_data = 12'b110011110111;
		14'b00101011001100: color_data = 12'b110011110111;
		14'b00101011001101: color_data = 12'b110011110111;
		14'b00101011001110: color_data = 12'b110011110111;
		14'b00101011001111: color_data = 12'b110011110111;
		14'b00101011010000: color_data = 12'b110011110111;
		14'b00101011010001: color_data = 12'b110011110111;
		14'b00101100000000: color_data = 12'b110011110111;
		14'b00101100000001: color_data = 12'b110011110111;
		14'b00101100000010: color_data = 12'b110011110111;
		14'b00101100000011: color_data = 12'b110011110111;
		14'b00101100000100: color_data = 12'b110011110111;
		14'b00101100000101: color_data = 12'b110011110111;
		14'b00101100001011: color_data = 12'b110011110111;
		14'b00101100001100: color_data = 12'b110011110111;
		14'b00101100001101: color_data = 12'b110011110111;
		14'b00101100001110: color_data = 12'b110011110111;
		14'b00101100001111: color_data = 12'b110011110111;
		14'b00101100010000: color_data = 12'b110011110111;
		14'b00101100010110: color_data = 12'b110011110111;
		14'b00101100010111: color_data = 12'b110011110111;
		14'b00101100011000: color_data = 12'b110011110111;
		14'b00101100011001: color_data = 12'b110011110111;
		14'b00101100011010: color_data = 12'b110011110111;
		14'b00101100100001: color_data = 12'b110011110111;
		14'b00101100100010: color_data = 12'b110011110111;
		14'b00101100100011: color_data = 12'b110011110111;
		14'b00101100100100: color_data = 12'b110011110111;
		14'b00101100100101: color_data = 12'b110011110111;
		14'b00101100101100: color_data = 12'b110011110111;
		14'b00101100101101: color_data = 12'b110011110111;
		14'b00101100101110: color_data = 12'b110011110111;
		14'b00101100101111: color_data = 12'b110011110111;
		14'b00101100110000: color_data = 12'b110011110111;
		14'b00101100110110: color_data = 12'b110011110111;
		14'b00101100110111: color_data = 12'b110011110111;
		14'b00101100111000: color_data = 12'b110011110111;
		14'b00101100111001: color_data = 12'b110011110111;
		14'b00101100111010: color_data = 12'b110011110111;
		14'b00101100111011: color_data = 12'b110011110111;
		14'b00101101000001: color_data = 12'b110011110111;
		14'b00101101000010: color_data = 12'b110011110111;
		14'b00101101000011: color_data = 12'b110011110111;
		14'b00101101000100: color_data = 12'b110011110111;
		14'b00101101000101: color_data = 12'b110011110111;
		14'b00101101000110: color_data = 12'b110011110111;
		14'b00101101000111: color_data = 12'b110011110111;
		14'b00101101001000: color_data = 12'b110011110111;
		14'b00101101001001: color_data = 12'b110011110111;
		14'b00101101001010: color_data = 12'b110011110111;
		14'b00101101001011: color_data = 12'b110011110111;
		14'b00101101010001: color_data = 12'b110011110111;
		14'b00101101010010: color_data = 12'b110011110111;
		14'b00101101010011: color_data = 12'b110011110111;
		14'b00101101010100: color_data = 12'b110011110111;
		14'b00101101010101: color_data = 12'b110011110111;
		14'b00101101010110: color_data = 12'b110011110111;
		14'b00101101100001: color_data = 12'b110011110111;
		14'b00101101100010: color_data = 12'b110011110111;
		14'b00101101100011: color_data = 12'b110011110111;
		14'b00101101100100: color_data = 12'b110011110111;
		14'b00101101100101: color_data = 12'b110011110111;
		14'b00101101100110: color_data = 12'b110011110111;
		14'b00101101100111: color_data = 12'b110011110111;
		14'b00101101101000: color_data = 12'b110011110111;
		14'b00101101101001: color_data = 12'b110011110111;
		14'b00101101101010: color_data = 12'b110011110111;
		14'b00101101101011: color_data = 12'b110011110111;
		14'b00101101101100: color_data = 12'b110011110111;
		14'b00101101101101: color_data = 12'b110011110111;
		14'b00101101101110: color_data = 12'b110011110111;
		14'b00101101101111: color_data = 12'b110011110111;
		14'b00101101110000: color_data = 12'b110011110111;
		14'b00101101110001: color_data = 12'b110011110111;
		14'b00101101110010: color_data = 12'b110011110111;
		14'b00101101110011: color_data = 12'b110011110111;
		14'b00101101110100: color_data = 12'b110011110111;
		14'b00101101110101: color_data = 12'b110011110111;
		14'b00101101110110: color_data = 12'b110011110111;
		14'b00101101111100: color_data = 12'b110011110111;
		14'b00101101111101: color_data = 12'b110011110111;
		14'b00101101111110: color_data = 12'b110011110111;
		14'b00101101111111: color_data = 12'b110011110111;
		14'b00101110000000: color_data = 12'b110011110111;
		14'b00101110000001: color_data = 12'b110011110111;
		14'b00101110001100: color_data = 12'b110011110111;
		14'b00101110001101: color_data = 12'b110011110111;
		14'b00101110001110: color_data = 12'b110011110111;
		14'b00101110001111: color_data = 12'b110011110111;
		14'b00101110010000: color_data = 12'b110011110111;
		14'b00101110010001: color_data = 12'b110011110111;
		14'b00101110010010: color_data = 12'b110011110111;
		14'b00101110010011: color_data = 12'b110011110111;
		14'b00101110010100: color_data = 12'b110011110111;
		14'b00101110010101: color_data = 12'b110011110111;
		14'b00101110010110: color_data = 12'b110011110111;
		14'b00101110011101: color_data = 12'b110011110111;
		14'b00101110011110: color_data = 12'b110011110111;
		14'b00101110011111: color_data = 12'b110011110111;
		14'b00101110100000: color_data = 12'b110011110111;
		14'b00101110100001: color_data = 12'b110011110111;
		14'b00101110100111: color_data = 12'b110011110111;
		14'b00101110101000: color_data = 12'b110011110111;
		14'b00101110101001: color_data = 12'b110011110111;
		14'b00101110101010: color_data = 12'b110011110111;
		14'b00101110101011: color_data = 12'b110011110111;
		14'b00101110101100: color_data = 12'b110011110111;
		14'b00101110110010: color_data = 12'b110011110111;
		14'b00101110110011: color_data = 12'b110011110111;
		14'b00101110110100: color_data = 12'b110011110111;
		14'b00101110110101: color_data = 12'b110011110111;
		14'b00101110110110: color_data = 12'b110011110111;
		14'b00101110110111: color_data = 12'b110011110111;
		14'b00101110111000: color_data = 12'b110011110111;
		14'b00101110111001: color_data = 12'b110011110111;
		14'b00101110111010: color_data = 12'b110011110111;
		14'b00101110111011: color_data = 12'b110011110111;
		14'b00101110111100: color_data = 12'b110011110111;
		14'b00101110111101: color_data = 12'b110011110111;
		14'b00101110111110: color_data = 12'b110011110111;
		14'b00101110111111: color_data = 12'b110011110111;
		14'b00101111000000: color_data = 12'b110011110111;
		14'b00101111000001: color_data = 12'b110011110111;
		14'b00101111001000: color_data = 12'b110011110111;
		14'b00101111001001: color_data = 12'b110011110111;
		14'b00101111001010: color_data = 12'b110011110111;
		14'b00101111001011: color_data = 12'b110011110111;
		14'b00101111001100: color_data = 12'b110011110111;
		14'b00101111001101: color_data = 12'b110011110111;
		14'b00101111001110: color_data = 12'b110011110111;
		14'b00101111001111: color_data = 12'b110011110111;
		14'b00101111010000: color_data = 12'b110011110111;
		14'b00101111010001: color_data = 12'b110011110111;
		14'b00110000000000: color_data = 12'b110011110111;
		14'b00110000000001: color_data = 12'b110011110111;
		14'b00110000000010: color_data = 12'b110011110111;
		14'b00110000000011: color_data = 12'b110011110111;
		14'b00110000000100: color_data = 12'b110011110111;
		14'b00110000000101: color_data = 12'b110011110111;
		14'b00110000001011: color_data = 12'b110011110111;
		14'b00110000001100: color_data = 12'b110011110111;
		14'b00110000001101: color_data = 12'b110011110111;
		14'b00110000001110: color_data = 12'b110011110111;
		14'b00110000001111: color_data = 12'b110011110111;
		14'b00110000010000: color_data = 12'b110011110111;
		14'b00110000010110: color_data = 12'b110011110111;
		14'b00110000010111: color_data = 12'b110011110111;
		14'b00110000011000: color_data = 12'b110011110111;
		14'b00110000011001: color_data = 12'b110011110111;
		14'b00110000011010: color_data = 12'b110011110111;
		14'b00110000100001: color_data = 12'b110011110111;
		14'b00110000100010: color_data = 12'b110011110111;
		14'b00110000100011: color_data = 12'b110011110111;
		14'b00110000100100: color_data = 12'b110011110111;
		14'b00110000100101: color_data = 12'b110011110111;
		14'b00110000101100: color_data = 12'b110011110111;
		14'b00110000101101: color_data = 12'b110011110111;
		14'b00110000101110: color_data = 12'b110011110111;
		14'b00110000101111: color_data = 12'b110011110111;
		14'b00110000110000: color_data = 12'b110011110111;
		14'b00110000110110: color_data = 12'b110011110111;
		14'b00110000110111: color_data = 12'b110011110111;
		14'b00110000111000: color_data = 12'b110011110111;
		14'b00110000111001: color_data = 12'b110011110111;
		14'b00110000111010: color_data = 12'b110011110111;
		14'b00110000111011: color_data = 12'b110011110111;
		14'b00110001000001: color_data = 12'b110011110111;
		14'b00110001000010: color_data = 12'b110011110111;
		14'b00110001000011: color_data = 12'b110011110111;
		14'b00110001000100: color_data = 12'b110011110111;
		14'b00110001000101: color_data = 12'b110011110111;
		14'b00110001000110: color_data = 12'b110011110111;
		14'b00110001000111: color_data = 12'b110011110111;
		14'b00110001001000: color_data = 12'b110011110111;
		14'b00110001001001: color_data = 12'b110011110111;
		14'b00110001001010: color_data = 12'b110011110111;
		14'b00110001001011: color_data = 12'b110011110111;
		14'b00110001010001: color_data = 12'b110011110111;
		14'b00110001010010: color_data = 12'b110011110111;
		14'b00110001010011: color_data = 12'b110011110111;
		14'b00110001010100: color_data = 12'b110011110111;
		14'b00110001010101: color_data = 12'b110011110111;
		14'b00110001010110: color_data = 12'b110011110111;
		14'b00110001100001: color_data = 12'b110011110111;
		14'b00110001100010: color_data = 12'b110011110111;
		14'b00110001100011: color_data = 12'b110011110111;
		14'b00110001100100: color_data = 12'b110011110111;
		14'b00110001100101: color_data = 12'b110011110111;
		14'b00110001100110: color_data = 12'b110011110111;
		14'b00110001100111: color_data = 12'b110011110111;
		14'b00110001101000: color_data = 12'b110011110111;
		14'b00110001101001: color_data = 12'b110011110111;
		14'b00110001101010: color_data = 12'b110011110111;
		14'b00110001101011: color_data = 12'b110011110111;
		14'b00110001101100: color_data = 12'b110011110111;
		14'b00110001101101: color_data = 12'b110011110111;
		14'b00110001101110: color_data = 12'b110011110111;
		14'b00110001101111: color_data = 12'b110011110111;
		14'b00110001110000: color_data = 12'b110011110111;
		14'b00110001110001: color_data = 12'b110011110111;
		14'b00110001110010: color_data = 12'b110011110111;
		14'b00110001110011: color_data = 12'b110011110111;
		14'b00110001110100: color_data = 12'b110011110111;
		14'b00110001110101: color_data = 12'b110011110111;
		14'b00110001110110: color_data = 12'b110011110111;
		14'b00110001111100: color_data = 12'b110011110111;
		14'b00110001111101: color_data = 12'b110011110111;
		14'b00110001111110: color_data = 12'b110011110111;
		14'b00110001111111: color_data = 12'b110011110111;
		14'b00110010000000: color_data = 12'b110011110111;
		14'b00110010000001: color_data = 12'b110011110111;
		14'b00110010001100: color_data = 12'b110011110111;
		14'b00110010001101: color_data = 12'b110011110111;
		14'b00110010001110: color_data = 12'b110011110111;
		14'b00110010001111: color_data = 12'b110011110111;
		14'b00110010010000: color_data = 12'b110011110111;
		14'b00110010010001: color_data = 12'b110011110111;
		14'b00110010010010: color_data = 12'b110011110111;
		14'b00110010010011: color_data = 12'b110011110111;
		14'b00110010010100: color_data = 12'b110011110111;
		14'b00110010010101: color_data = 12'b110011110111;
		14'b00110010010110: color_data = 12'b110011110111;
		14'b00110010011101: color_data = 12'b110011110111;
		14'b00110010011110: color_data = 12'b110011110111;
		14'b00110010011111: color_data = 12'b110011110111;
		14'b00110010100000: color_data = 12'b110011110111;
		14'b00110010100001: color_data = 12'b110011110111;
		14'b00110010100111: color_data = 12'b110011110111;
		14'b00110010101000: color_data = 12'b110011110111;
		14'b00110010101001: color_data = 12'b110011110111;
		14'b00110010101010: color_data = 12'b110011110111;
		14'b00110010101011: color_data = 12'b110011110111;
		14'b00110010101100: color_data = 12'b110011110111;
		14'b00110010110010: color_data = 12'b110011110111;
		14'b00110010110011: color_data = 12'b110011110111;
		14'b00110010110100: color_data = 12'b110011110111;
		14'b00110010110101: color_data = 12'b110011110111;
		14'b00110010110110: color_data = 12'b110011110111;
		14'b00110010110111: color_data = 12'b110011110111;
		14'b00110010111000: color_data = 12'b110011110111;
		14'b00110010111001: color_data = 12'b110011110111;
		14'b00110010111010: color_data = 12'b110011110111;
		14'b00110010111011: color_data = 12'b110011110111;
		14'b00110010111100: color_data = 12'b110011110111;
		14'b00110010111101: color_data = 12'b110011110111;
		14'b00110010111110: color_data = 12'b110011110111;
		14'b00110010111111: color_data = 12'b110011110111;
		14'b00110011000000: color_data = 12'b110011110111;
		14'b00110011000001: color_data = 12'b110011110111;
		14'b00110011001000: color_data = 12'b110011110111;
		14'b00110011001001: color_data = 12'b110011110111;
		14'b00110011001010: color_data = 12'b110011110111;
		14'b00110011001011: color_data = 12'b110011110111;
		14'b00110011001100: color_data = 12'b110011110111;
		14'b00110011001101: color_data = 12'b110011110111;
		14'b00110011001110: color_data = 12'b110011110111;
		14'b00110011001111: color_data = 12'b110011110111;
		14'b00110011010000: color_data = 12'b110011110111;
		14'b00110011010001: color_data = 12'b110011110111;
		14'b00110100000000: color_data = 12'b110011110111;
		14'b00110100000001: color_data = 12'b110011110111;
		14'b00110100000010: color_data = 12'b110011110111;
		14'b00110100000011: color_data = 12'b110011110111;
		14'b00110100000100: color_data = 12'b110011110111;
		14'b00110100000101: color_data = 12'b110011110111;
		14'b00110100001011: color_data = 12'b110011110111;
		14'b00110100001100: color_data = 12'b110011110111;
		14'b00110100001101: color_data = 12'b110011110111;
		14'b00110100001110: color_data = 12'b110011110111;
		14'b00110100001111: color_data = 12'b110011110111;
		14'b00110100010000: color_data = 12'b110011110111;
		14'b00110100010110: color_data = 12'b110011110111;
		14'b00110100010111: color_data = 12'b110011110111;
		14'b00110100011000: color_data = 12'b110011110111;
		14'b00110100011001: color_data = 12'b110011110111;
		14'b00110100011010: color_data = 12'b110011110111;
		14'b00110100100001: color_data = 12'b110011110111;
		14'b00110100100010: color_data = 12'b110011110111;
		14'b00110100100011: color_data = 12'b110011110111;
		14'b00110100100100: color_data = 12'b110011110111;
		14'b00110100100101: color_data = 12'b110011110111;
		14'b00110100101100: color_data = 12'b110011110111;
		14'b00110100101101: color_data = 12'b110011110111;
		14'b00110100101110: color_data = 12'b110011110111;
		14'b00110100101111: color_data = 12'b110011110111;
		14'b00110100110000: color_data = 12'b110011110111;
		14'b00110100110110: color_data = 12'b110011110111;
		14'b00110100110111: color_data = 12'b110011110111;
		14'b00110100111000: color_data = 12'b110011110111;
		14'b00110100111001: color_data = 12'b110011110111;
		14'b00110100111010: color_data = 12'b110011110111;
		14'b00110100111011: color_data = 12'b110011110111;
		14'b00110101000001: color_data = 12'b110011110111;
		14'b00110101000010: color_data = 12'b110011110111;
		14'b00110101000011: color_data = 12'b110011110111;
		14'b00110101000100: color_data = 12'b110011110111;
		14'b00110101000101: color_data = 12'b110011110111;
		14'b00110101000110: color_data = 12'b110011110111;
		14'b00110101000111: color_data = 12'b110011110111;
		14'b00110101001000: color_data = 12'b110011110111;
		14'b00110101001001: color_data = 12'b110011110111;
		14'b00110101001010: color_data = 12'b110011110111;
		14'b00110101001011: color_data = 12'b110011110111;
		14'b00110101010001: color_data = 12'b110011110111;
		14'b00110101010010: color_data = 12'b110011110111;
		14'b00110101010011: color_data = 12'b110011110111;
		14'b00110101010100: color_data = 12'b110011110111;
		14'b00110101010101: color_data = 12'b110011110111;
		14'b00110101010110: color_data = 12'b110011110111;
		14'b00110101100001: color_data = 12'b110011110111;
		14'b00110101100010: color_data = 12'b110011110111;
		14'b00110101100011: color_data = 12'b110011110111;
		14'b00110101100100: color_data = 12'b110011110111;
		14'b00110101100101: color_data = 12'b110011110111;
		14'b00110101100110: color_data = 12'b110011110111;
		14'b00110101100111: color_data = 12'b110011110111;
		14'b00110101101000: color_data = 12'b110011110111;
		14'b00110101101001: color_data = 12'b110011110111;
		14'b00110101101010: color_data = 12'b110011110111;
		14'b00110101101011: color_data = 12'b110011110111;
		14'b00110101101100: color_data = 12'b110011110111;
		14'b00110101101101: color_data = 12'b110011110111;
		14'b00110101101110: color_data = 12'b110011110111;
		14'b00110101101111: color_data = 12'b110011110111;
		14'b00110101110000: color_data = 12'b110011110111;
		14'b00110101110001: color_data = 12'b110011110111;
		14'b00110101110010: color_data = 12'b110011110111;
		14'b00110101110011: color_data = 12'b110011110111;
		14'b00110101110100: color_data = 12'b110011110111;
		14'b00110101110101: color_data = 12'b110011110111;
		14'b00110101110110: color_data = 12'b110011110111;
		14'b00110101111100: color_data = 12'b110011110111;
		14'b00110101111101: color_data = 12'b110011110111;
		14'b00110101111110: color_data = 12'b110011110111;
		14'b00110101111111: color_data = 12'b110011110111;
		14'b00110110000000: color_data = 12'b110011110111;
		14'b00110110000001: color_data = 12'b110011110111;
		14'b00110110001100: color_data = 12'b110011110111;
		14'b00110110001101: color_data = 12'b110011110111;
		14'b00110110001110: color_data = 12'b110011110111;
		14'b00110110001111: color_data = 12'b110011110111;
		14'b00110110010000: color_data = 12'b110011110111;
		14'b00110110010001: color_data = 12'b110011110111;
		14'b00110110010010: color_data = 12'b110011110111;
		14'b00110110010011: color_data = 12'b110011110111;
		14'b00110110010100: color_data = 12'b110011110111;
		14'b00110110010101: color_data = 12'b110011110111;
		14'b00110110010110: color_data = 12'b110011110111;
		14'b00110110011101: color_data = 12'b110011110111;
		14'b00110110011110: color_data = 12'b110011110111;
		14'b00110110011111: color_data = 12'b110011110111;
		14'b00110110100000: color_data = 12'b110011110111;
		14'b00110110100001: color_data = 12'b110011110111;
		14'b00110110100111: color_data = 12'b110011110111;
		14'b00110110101000: color_data = 12'b110011110111;
		14'b00110110101001: color_data = 12'b110011110111;
		14'b00110110101010: color_data = 12'b110011110111;
		14'b00110110101011: color_data = 12'b110011110111;
		14'b00110110101100: color_data = 12'b110011110111;
		14'b00110110110010: color_data = 12'b110011110111;
		14'b00110110110011: color_data = 12'b110011110111;
		14'b00110110110100: color_data = 12'b110011110111;
		14'b00110110110101: color_data = 12'b110011110111;
		14'b00110110110110: color_data = 12'b110011110111;
		14'b00110110110111: color_data = 12'b110011110111;
		14'b00110110111000: color_data = 12'b110011110111;
		14'b00110110111001: color_data = 12'b110011110111;
		14'b00110110111010: color_data = 12'b110011110111;
		14'b00110110111011: color_data = 12'b110011110111;
		14'b00110110111100: color_data = 12'b110011110111;
		14'b00110110111101: color_data = 12'b110011110111;
		14'b00110110111110: color_data = 12'b110011110111;
		14'b00110110111111: color_data = 12'b110011110111;
		14'b00110111000000: color_data = 12'b110011110111;
		14'b00110111000001: color_data = 12'b110011110111;
		14'b00110111001000: color_data = 12'b110011110111;
		14'b00110111001001: color_data = 12'b110011110111;
		14'b00110111001010: color_data = 12'b110011110111;
		14'b00110111001011: color_data = 12'b110011110111;
		14'b00110111001100: color_data = 12'b110011110111;
		14'b00110111001101: color_data = 12'b110011110111;
		14'b00110111001110: color_data = 12'b110011110111;
		14'b00110111001111: color_data = 12'b110011110111;
		14'b00110111010000: color_data = 12'b110011110111;
		14'b00110111010001: color_data = 12'b110011110111;
		14'b00111000000000: color_data = 12'b110011110111;
		14'b00111000000001: color_data = 12'b110011110111;
		14'b00111000000010: color_data = 12'b110011110111;
		14'b00111000000011: color_data = 12'b110011110111;
		14'b00111000000100: color_data = 12'b110011110111;
		14'b00111000000101: color_data = 12'b110011110111;
		14'b00111000001011: color_data = 12'b110011110111;
		14'b00111000001100: color_data = 12'b110011110111;
		14'b00111000001101: color_data = 12'b110011110111;
		14'b00111000001110: color_data = 12'b110011110111;
		14'b00111000001111: color_data = 12'b110011110111;
		14'b00111000010000: color_data = 12'b110011110111;
		14'b00111000010110: color_data = 12'b110011110111;
		14'b00111000010111: color_data = 12'b110011110111;
		14'b00111000011000: color_data = 12'b110011110111;
		14'b00111000011001: color_data = 12'b110011110111;
		14'b00111000011010: color_data = 12'b110011110111;
		14'b00111000100001: color_data = 12'b110011110111;
		14'b00111000100010: color_data = 12'b110011110111;
		14'b00111000100011: color_data = 12'b110011110111;
		14'b00111000100100: color_data = 12'b110011110111;
		14'b00111000100101: color_data = 12'b110011110111;
		14'b00111000101100: color_data = 12'b110011110111;
		14'b00111000101101: color_data = 12'b110011110111;
		14'b00111000101110: color_data = 12'b110011110111;
		14'b00111000101111: color_data = 12'b110011110111;
		14'b00111000110000: color_data = 12'b110011110111;
		14'b00111000110110: color_data = 12'b110011110111;
		14'b00111000110111: color_data = 12'b110011110111;
		14'b00111000111000: color_data = 12'b110011110111;
		14'b00111000111001: color_data = 12'b110011110111;
		14'b00111000111010: color_data = 12'b110011110111;
		14'b00111000111011: color_data = 12'b110011110111;
		14'b00111001000001: color_data = 12'b110011110111;
		14'b00111001000010: color_data = 12'b110011110111;
		14'b00111001000011: color_data = 12'b110011110111;
		14'b00111001000100: color_data = 12'b110011110111;
		14'b00111001000101: color_data = 12'b110011110111;
		14'b00111001010001: color_data = 12'b110011110111;
		14'b00111001010010: color_data = 12'b110011110111;
		14'b00111001010011: color_data = 12'b110011110111;
		14'b00111001010100: color_data = 12'b110011110111;
		14'b00111001010101: color_data = 12'b110011110111;
		14'b00111001010110: color_data = 12'b110011110111;
		14'b00111001100001: color_data = 12'b110011110111;
		14'b00111001100010: color_data = 12'b110011110111;
		14'b00111001100011: color_data = 12'b110011110111;
		14'b00111001100100: color_data = 12'b110011110111;
		14'b00111001100101: color_data = 12'b110011110111;
		14'b00111001100110: color_data = 12'b110011110111;
		14'b00111001111100: color_data = 12'b110011110111;
		14'b00111001111101: color_data = 12'b110011110111;
		14'b00111001111110: color_data = 12'b110011110111;
		14'b00111001111111: color_data = 12'b110011110111;
		14'b00111010000000: color_data = 12'b110011110111;
		14'b00111010000001: color_data = 12'b110011110111;
		14'b00111010000111: color_data = 12'b110011110111;
		14'b00111010001000: color_data = 12'b110011110111;
		14'b00111010001001: color_data = 12'b110011110111;
		14'b00111010001010: color_data = 12'b110011110111;
		14'b00111010001011: color_data = 12'b110011110111;
		14'b00111010010010: color_data = 12'b110011110111;
		14'b00111010010011: color_data = 12'b110011110111;
		14'b00111010010100: color_data = 12'b110011110111;
		14'b00111010010101: color_data = 12'b110011110111;
		14'b00111010010110: color_data = 12'b110011110111;
		14'b00111010011101: color_data = 12'b110011110111;
		14'b00111010011110: color_data = 12'b110011110111;
		14'b00111010011111: color_data = 12'b110011110111;
		14'b00111010100000: color_data = 12'b110011110111;
		14'b00111010100001: color_data = 12'b110011110111;
		14'b00111010100111: color_data = 12'b110011110111;
		14'b00111010101000: color_data = 12'b110011110111;
		14'b00111010101001: color_data = 12'b110011110111;
		14'b00111010101010: color_data = 12'b110011110111;
		14'b00111010101011: color_data = 12'b110011110111;
		14'b00111010101100: color_data = 12'b110011110111;
		14'b00111010110010: color_data = 12'b110011110111;
		14'b00111010110011: color_data = 12'b110011110111;
		14'b00111010110100: color_data = 12'b110011110111;
		14'b00111010110101: color_data = 12'b110011110111;
		14'b00111010110110: color_data = 12'b110011110111;
		14'b00111010110111: color_data = 12'b110011110111;
		14'b00111010111101: color_data = 12'b110011110111;
		14'b00111010111110: color_data = 12'b110011110111;
		14'b00111010111111: color_data = 12'b110011110111;
		14'b00111011000000: color_data = 12'b110011110111;
		14'b00111011000001: color_data = 12'b110011110111;
		14'b00111011001000: color_data = 12'b110011110111;
		14'b00111011001001: color_data = 12'b110011110111;
		14'b00111011001010: color_data = 12'b110011110111;
		14'b00111011001011: color_data = 12'b110011110111;
		14'b00111011001100: color_data = 12'b110011110111;
		14'b00111100000000: color_data = 12'b110011110111;
		14'b00111100000001: color_data = 12'b110011110111;
		14'b00111100000010: color_data = 12'b110011110111;
		14'b00111100000011: color_data = 12'b110011110111;
		14'b00111100000100: color_data = 12'b110011110111;
		14'b00111100000101: color_data = 12'b110011110111;
		14'b00111100001011: color_data = 12'b110011110111;
		14'b00111100001100: color_data = 12'b110011110111;
		14'b00111100001101: color_data = 12'b110011110111;
		14'b00111100001110: color_data = 12'b110011110111;
		14'b00111100001111: color_data = 12'b110011110111;
		14'b00111100010000: color_data = 12'b110011110111;
		14'b00111100010110: color_data = 12'b110011110111;
		14'b00111100010111: color_data = 12'b110011110111;
		14'b00111100011000: color_data = 12'b110011110111;
		14'b00111100011001: color_data = 12'b110011110111;
		14'b00111100011010: color_data = 12'b110011110111;
		14'b00111100100001: color_data = 12'b110011110111;
		14'b00111100100010: color_data = 12'b110011110111;
		14'b00111100100011: color_data = 12'b110011110111;
		14'b00111100100100: color_data = 12'b110011110111;
		14'b00111100100101: color_data = 12'b110011110111;
		14'b00111100101100: color_data = 12'b110011110111;
		14'b00111100101101: color_data = 12'b110011110111;
		14'b00111100101110: color_data = 12'b110011110111;
		14'b00111100101111: color_data = 12'b110011110111;
		14'b00111100110000: color_data = 12'b110011110111;
		14'b00111100110110: color_data = 12'b110011110111;
		14'b00111100110111: color_data = 12'b110011110111;
		14'b00111100111000: color_data = 12'b110011110111;
		14'b00111100111001: color_data = 12'b110011110111;
		14'b00111100111010: color_data = 12'b110011110111;
		14'b00111100111011: color_data = 12'b110011110111;
		14'b00111101000001: color_data = 12'b110011110111;
		14'b00111101000010: color_data = 12'b110011110111;
		14'b00111101000011: color_data = 12'b110011110111;
		14'b00111101000100: color_data = 12'b110011110111;
		14'b00111101000101: color_data = 12'b110011110111;
		14'b00111101010001: color_data = 12'b110011110111;
		14'b00111101010010: color_data = 12'b110011110111;
		14'b00111101010011: color_data = 12'b110011110111;
		14'b00111101010100: color_data = 12'b110011110111;
		14'b00111101010101: color_data = 12'b110011110111;
		14'b00111101010110: color_data = 12'b110011110111;
		14'b00111101100001: color_data = 12'b110011110111;
		14'b00111101100010: color_data = 12'b110011110111;
		14'b00111101100011: color_data = 12'b110011110111;
		14'b00111101100100: color_data = 12'b110011110111;
		14'b00111101100101: color_data = 12'b110011110111;
		14'b00111101100110: color_data = 12'b110011110111;
		14'b00111101111100: color_data = 12'b110011110111;
		14'b00111101111101: color_data = 12'b110011110111;
		14'b00111101111110: color_data = 12'b110011110111;
		14'b00111101111111: color_data = 12'b110011110111;
		14'b00111110000000: color_data = 12'b110011110111;
		14'b00111110000001: color_data = 12'b110011110111;
		14'b00111110000111: color_data = 12'b110011110111;
		14'b00111110001000: color_data = 12'b110011110111;
		14'b00111110001001: color_data = 12'b110011110111;
		14'b00111110001010: color_data = 12'b110011110111;
		14'b00111110001011: color_data = 12'b110011110111;
		14'b00111110010010: color_data = 12'b110011110111;
		14'b00111110010011: color_data = 12'b110011110111;
		14'b00111110010100: color_data = 12'b110011110111;
		14'b00111110010101: color_data = 12'b110011110111;
		14'b00111110010110: color_data = 12'b110011110111;
		14'b00111110011101: color_data = 12'b110011110111;
		14'b00111110011110: color_data = 12'b110011110111;
		14'b00111110011111: color_data = 12'b110011110111;
		14'b00111110100000: color_data = 12'b110011110111;
		14'b00111110100001: color_data = 12'b110011110111;
		14'b00111110100111: color_data = 12'b110011110111;
		14'b00111110101000: color_data = 12'b110011110111;
		14'b00111110101001: color_data = 12'b110011110111;
		14'b00111110101010: color_data = 12'b110011110111;
		14'b00111110101011: color_data = 12'b110011110111;
		14'b00111110101100: color_data = 12'b110011110111;
		14'b00111110110010: color_data = 12'b110011110111;
		14'b00111110110011: color_data = 12'b110011110111;
		14'b00111110110100: color_data = 12'b110011110111;
		14'b00111110110101: color_data = 12'b110011110111;
		14'b00111110110110: color_data = 12'b110011110111;
		14'b00111110110111: color_data = 12'b110011110111;
		14'b00111110111101: color_data = 12'b110011110111;
		14'b00111110111110: color_data = 12'b110011110111;
		14'b00111110111111: color_data = 12'b110011110111;
		14'b00111111000000: color_data = 12'b110011110111;
		14'b00111111000001: color_data = 12'b110011110111;
		14'b00111111001000: color_data = 12'b110011110111;
		14'b00111111001001: color_data = 12'b110011110111;
		14'b00111111001010: color_data = 12'b110011110111;
		14'b00111111001011: color_data = 12'b110011110111;
		14'b00111111001100: color_data = 12'b110011110111;
		14'b01000000000000: color_data = 12'b110011110111;
		14'b01000000000001: color_data = 12'b110011110111;
		14'b01000000000010: color_data = 12'b110011110111;
		14'b01000000000011: color_data = 12'b110011110111;
		14'b01000000000100: color_data = 12'b110011110111;
		14'b01000000000101: color_data = 12'b110011110111;
		14'b01000000001011: color_data = 12'b110011110111;
		14'b01000000001100: color_data = 12'b110011110111;
		14'b01000000001101: color_data = 12'b110011110111;
		14'b01000000001110: color_data = 12'b110011110111;
		14'b01000000001111: color_data = 12'b110011110111;
		14'b01000000010000: color_data = 12'b110011110111;
		14'b01000000010110: color_data = 12'b110011110111;
		14'b01000000010111: color_data = 12'b110011110111;
		14'b01000000011000: color_data = 12'b110011110111;
		14'b01000000011001: color_data = 12'b110011110111;
		14'b01000000011010: color_data = 12'b110011110111;
		14'b01000000100001: color_data = 12'b110011110111;
		14'b01000000100010: color_data = 12'b110011110111;
		14'b01000000100011: color_data = 12'b110011110111;
		14'b01000000100100: color_data = 12'b110011110111;
		14'b01000000100101: color_data = 12'b110011110111;
		14'b01000000101100: color_data = 12'b110011110111;
		14'b01000000101101: color_data = 12'b110011110111;
		14'b01000000101110: color_data = 12'b110011110111;
		14'b01000000101111: color_data = 12'b110011110111;
		14'b01000000110000: color_data = 12'b110011110111;
		14'b01000000110110: color_data = 12'b110011110111;
		14'b01000000110111: color_data = 12'b110011110111;
		14'b01000000111000: color_data = 12'b110011110111;
		14'b01000000111001: color_data = 12'b110011110111;
		14'b01000000111010: color_data = 12'b110011110111;
		14'b01000000111011: color_data = 12'b110011110111;
		14'b01000001000001: color_data = 12'b110011110111;
		14'b01000001000010: color_data = 12'b110011110111;
		14'b01000001000011: color_data = 12'b110011110111;
		14'b01000001000100: color_data = 12'b110011110111;
		14'b01000001000101: color_data = 12'b110011110111;
		14'b01000001010001: color_data = 12'b110011110111;
		14'b01000001010010: color_data = 12'b110011110111;
		14'b01000001010011: color_data = 12'b110011110111;
		14'b01000001010100: color_data = 12'b110011110111;
		14'b01000001010101: color_data = 12'b110011110111;
		14'b01000001010110: color_data = 12'b110011110111;
		14'b01000001100001: color_data = 12'b110011110111;
		14'b01000001100010: color_data = 12'b110011110111;
		14'b01000001100011: color_data = 12'b110011110111;
		14'b01000001100100: color_data = 12'b110011110111;
		14'b01000001100101: color_data = 12'b110011110111;
		14'b01000001100110: color_data = 12'b110011110111;
		14'b01000001111100: color_data = 12'b110011110111;
		14'b01000001111101: color_data = 12'b110011110111;
		14'b01000001111110: color_data = 12'b110011110111;
		14'b01000001111111: color_data = 12'b110011110111;
		14'b01000010000000: color_data = 12'b110011110111;
		14'b01000010000001: color_data = 12'b110011110111;
		14'b01000010000111: color_data = 12'b110011110111;
		14'b01000010001000: color_data = 12'b110011110111;
		14'b01000010001001: color_data = 12'b110011110111;
		14'b01000010001010: color_data = 12'b110011110111;
		14'b01000010001011: color_data = 12'b110011110111;
		14'b01000010010010: color_data = 12'b110011110111;
		14'b01000010010011: color_data = 12'b110011110111;
		14'b01000010010100: color_data = 12'b110011110111;
		14'b01000010010101: color_data = 12'b110011110111;
		14'b01000010010110: color_data = 12'b110011110111;
		14'b01000010011101: color_data = 12'b110011110111;
		14'b01000010011110: color_data = 12'b110011110111;
		14'b01000010011111: color_data = 12'b110011110111;
		14'b01000010100000: color_data = 12'b110011110111;
		14'b01000010100001: color_data = 12'b110011110111;
		14'b01000010100111: color_data = 12'b110011110111;
		14'b01000010101000: color_data = 12'b110011110111;
		14'b01000010101001: color_data = 12'b110011110111;
		14'b01000010101010: color_data = 12'b110011110111;
		14'b01000010101011: color_data = 12'b110011110111;
		14'b01000010101100: color_data = 12'b110011110111;
		14'b01000010110010: color_data = 12'b110011110111;
		14'b01000010110011: color_data = 12'b110011110111;
		14'b01000010110100: color_data = 12'b110011110111;
		14'b01000010110101: color_data = 12'b110011110111;
		14'b01000010110110: color_data = 12'b110011110111;
		14'b01000010110111: color_data = 12'b110011110111;
		14'b01000010111101: color_data = 12'b110011110111;
		14'b01000010111110: color_data = 12'b110011110111;
		14'b01000010111111: color_data = 12'b110011110111;
		14'b01000011000000: color_data = 12'b110011110111;
		14'b01000011000001: color_data = 12'b110011110111;
		14'b01000011001000: color_data = 12'b110011110111;
		14'b01000011001001: color_data = 12'b110011110111;
		14'b01000011001010: color_data = 12'b110011110111;
		14'b01000011001011: color_data = 12'b110011110111;
		14'b01000011001100: color_data = 12'b110011110111;
		14'b01000100000000: color_data = 12'b110011110111;
		14'b01000100000001: color_data = 12'b110011110111;
		14'b01000100000010: color_data = 12'b110011110111;
		14'b01000100000011: color_data = 12'b110011110111;
		14'b01000100000100: color_data = 12'b110011110111;
		14'b01000100000101: color_data = 12'b110011110111;
		14'b01000100001011: color_data = 12'b110011110111;
		14'b01000100001100: color_data = 12'b110011110111;
		14'b01000100001101: color_data = 12'b110011110111;
		14'b01000100001110: color_data = 12'b110011110111;
		14'b01000100001111: color_data = 12'b110011110111;
		14'b01000100010000: color_data = 12'b110011110111;
		14'b01000100010110: color_data = 12'b110011110111;
		14'b01000100010111: color_data = 12'b110011110111;
		14'b01000100011000: color_data = 12'b110011110111;
		14'b01000100011001: color_data = 12'b110011110111;
		14'b01000100011010: color_data = 12'b110011110111;
		14'b01000100100001: color_data = 12'b110011110111;
		14'b01000100100010: color_data = 12'b110011110111;
		14'b01000100100011: color_data = 12'b110011110111;
		14'b01000100100100: color_data = 12'b110011110111;
		14'b01000100100101: color_data = 12'b110011110111;
		14'b01000100101100: color_data = 12'b110011110111;
		14'b01000100101101: color_data = 12'b110011110111;
		14'b01000100101110: color_data = 12'b110011110111;
		14'b01000100101111: color_data = 12'b110011110111;
		14'b01000100110000: color_data = 12'b110011110111;
		14'b01000100110110: color_data = 12'b110011110111;
		14'b01000100110111: color_data = 12'b110011110111;
		14'b01000100111000: color_data = 12'b110011110111;
		14'b01000100111001: color_data = 12'b110011110111;
		14'b01000100111010: color_data = 12'b110011110111;
		14'b01000100111011: color_data = 12'b110011110111;
		14'b01000101000001: color_data = 12'b110011110111;
		14'b01000101000010: color_data = 12'b110011110111;
		14'b01000101000011: color_data = 12'b110011110111;
		14'b01000101000100: color_data = 12'b110011110111;
		14'b01000101000101: color_data = 12'b110011110111;
		14'b01000101010001: color_data = 12'b110011110111;
		14'b01000101010010: color_data = 12'b110011110111;
		14'b01000101010011: color_data = 12'b110011110111;
		14'b01000101010100: color_data = 12'b110011110111;
		14'b01000101010101: color_data = 12'b110011110111;
		14'b01000101010110: color_data = 12'b110011110111;
		14'b01000101100001: color_data = 12'b110011110111;
		14'b01000101100010: color_data = 12'b110011110111;
		14'b01000101100011: color_data = 12'b110011110111;
		14'b01000101100100: color_data = 12'b110011110111;
		14'b01000101100101: color_data = 12'b110011110111;
		14'b01000101100110: color_data = 12'b110011110111;
		14'b01000101111100: color_data = 12'b110011110111;
		14'b01000101111101: color_data = 12'b110011110111;
		14'b01000101111110: color_data = 12'b110011110111;
		14'b01000101111111: color_data = 12'b110011110111;
		14'b01000110000000: color_data = 12'b110011110111;
		14'b01000110000001: color_data = 12'b110011110111;
		14'b01000110000111: color_data = 12'b110011110111;
		14'b01000110001000: color_data = 12'b110011110111;
		14'b01000110001001: color_data = 12'b110011110111;
		14'b01000110001010: color_data = 12'b110011110111;
		14'b01000110001011: color_data = 12'b110011110111;
		14'b01000110010010: color_data = 12'b110011110111;
		14'b01000110010011: color_data = 12'b110011110111;
		14'b01000110010100: color_data = 12'b110011110111;
		14'b01000110010101: color_data = 12'b110011110111;
		14'b01000110010110: color_data = 12'b110011110111;
		14'b01000110011101: color_data = 12'b110011110111;
		14'b01000110011110: color_data = 12'b110011110111;
		14'b01000110011111: color_data = 12'b110011110111;
		14'b01000110100000: color_data = 12'b110011110111;
		14'b01000110100001: color_data = 12'b110011110111;
		14'b01000110100111: color_data = 12'b110011110111;
		14'b01000110101000: color_data = 12'b110011110111;
		14'b01000110101001: color_data = 12'b110011110111;
		14'b01000110101010: color_data = 12'b110011110111;
		14'b01000110101011: color_data = 12'b110011110111;
		14'b01000110101100: color_data = 12'b110011110111;
		14'b01000110110010: color_data = 12'b110011110111;
		14'b01000110110011: color_data = 12'b110011110111;
		14'b01000110110100: color_data = 12'b110011110111;
		14'b01000110110101: color_data = 12'b110011110111;
		14'b01000110110110: color_data = 12'b110011110111;
		14'b01000110110111: color_data = 12'b110011110111;
		14'b01000110111101: color_data = 12'b110011110111;
		14'b01000110111110: color_data = 12'b110011110111;
		14'b01000110111111: color_data = 12'b110011110111;
		14'b01000111000000: color_data = 12'b110011110111;
		14'b01000111000001: color_data = 12'b110011110111;
		14'b01000111001000: color_data = 12'b110011110111;
		14'b01000111001001: color_data = 12'b110011110111;
		14'b01000111001010: color_data = 12'b110011110111;
		14'b01000111001011: color_data = 12'b110011110111;
		14'b01000111001100: color_data = 12'b110011110111;
		14'b01001000000000: color_data = 12'b110011110111;
		14'b01001000000001: color_data = 12'b110011110111;
		14'b01001000000010: color_data = 12'b110011110111;
		14'b01001000000011: color_data = 12'b110011110111;
		14'b01001000000100: color_data = 12'b110011110111;
		14'b01001000000101: color_data = 12'b110011110111;
		14'b01001000001011: color_data = 12'b110011110111;
		14'b01001000001100: color_data = 12'b110011110111;
		14'b01001000001101: color_data = 12'b110011110111;
		14'b01001000001110: color_data = 12'b110011110111;
		14'b01001000001111: color_data = 12'b110011110111;
		14'b01001000010000: color_data = 12'b110011110111;
		14'b01001000010110: color_data = 12'b110011110111;
		14'b01001000010111: color_data = 12'b110011110111;
		14'b01001000011000: color_data = 12'b110011110111;
		14'b01001000011001: color_data = 12'b110011110111;
		14'b01001000011010: color_data = 12'b110011110111;
		14'b01001000100001: color_data = 12'b110011110111;
		14'b01001000100010: color_data = 12'b110011110111;
		14'b01001000100011: color_data = 12'b110011110111;
		14'b01001000100100: color_data = 12'b110011110111;
		14'b01001000100101: color_data = 12'b110011110111;
		14'b01001000101100: color_data = 12'b110011110111;
		14'b01001000101101: color_data = 12'b110011110111;
		14'b01001000101110: color_data = 12'b110011110111;
		14'b01001000101111: color_data = 12'b110011110111;
		14'b01001000110000: color_data = 12'b110011110111;
		14'b01001000110110: color_data = 12'b110011110111;
		14'b01001000110111: color_data = 12'b110011110111;
		14'b01001000111000: color_data = 12'b110011110111;
		14'b01001000111001: color_data = 12'b110011110111;
		14'b01001000111010: color_data = 12'b110011110111;
		14'b01001000111011: color_data = 12'b110011110111;
		14'b01001001000001: color_data = 12'b110011110111;
		14'b01001001000010: color_data = 12'b110011110111;
		14'b01001001000011: color_data = 12'b110011110111;
		14'b01001001000100: color_data = 12'b110011110111;
		14'b01001001000101: color_data = 12'b110011110111;
		14'b01001001010001: color_data = 12'b110011110111;
		14'b01001001010010: color_data = 12'b110011110111;
		14'b01001001010011: color_data = 12'b110011110111;
		14'b01001001010100: color_data = 12'b110011110111;
		14'b01001001010101: color_data = 12'b110011110111;
		14'b01001001010110: color_data = 12'b110011110111;
		14'b01001001100001: color_data = 12'b110011110111;
		14'b01001001100010: color_data = 12'b110011110111;
		14'b01001001100011: color_data = 12'b110011110111;
		14'b01001001100100: color_data = 12'b110011110111;
		14'b01001001100101: color_data = 12'b110011110111;
		14'b01001001100110: color_data = 12'b110011110111;
		14'b01001001111100: color_data = 12'b110011110111;
		14'b01001001111101: color_data = 12'b110011110111;
		14'b01001001111110: color_data = 12'b110011110111;
		14'b01001001111111: color_data = 12'b110011110111;
		14'b01001010000000: color_data = 12'b110011110111;
		14'b01001010000001: color_data = 12'b110011110111;
		14'b01001010000111: color_data = 12'b110011110111;
		14'b01001010001000: color_data = 12'b110011110111;
		14'b01001010001001: color_data = 12'b110011110111;
		14'b01001010001010: color_data = 12'b110011110111;
		14'b01001010001011: color_data = 12'b110011110111;
		14'b01001010010010: color_data = 12'b110011110111;
		14'b01001010010011: color_data = 12'b110011110111;
		14'b01001010010100: color_data = 12'b110011110111;
		14'b01001010010101: color_data = 12'b110011110111;
		14'b01001010010110: color_data = 12'b110011110111;
		14'b01001010011101: color_data = 12'b110011110111;
		14'b01001010011110: color_data = 12'b110011110111;
		14'b01001010011111: color_data = 12'b110011110111;
		14'b01001010100000: color_data = 12'b110011110111;
		14'b01001010100001: color_data = 12'b110011110111;
		14'b01001010100111: color_data = 12'b110011110111;
		14'b01001010101000: color_data = 12'b110011110111;
		14'b01001010101001: color_data = 12'b110011110111;
		14'b01001010101010: color_data = 12'b110011110111;
		14'b01001010101011: color_data = 12'b110011110111;
		14'b01001010101100: color_data = 12'b110011110111;
		14'b01001010110010: color_data = 12'b110011110111;
		14'b01001010110011: color_data = 12'b110011110111;
		14'b01001010110100: color_data = 12'b110011110111;
		14'b01001010110101: color_data = 12'b110011110111;
		14'b01001010110110: color_data = 12'b110011110111;
		14'b01001010110111: color_data = 12'b110011110111;
		14'b01001010111101: color_data = 12'b110011110111;
		14'b01001010111110: color_data = 12'b110011110111;
		14'b01001010111111: color_data = 12'b110011110111;
		14'b01001011000000: color_data = 12'b110011110111;
		14'b01001011000001: color_data = 12'b110011110111;
		14'b01001011001000: color_data = 12'b110011110111;
		14'b01001011001001: color_data = 12'b110011110111;
		14'b01001011001010: color_data = 12'b110011110111;
		14'b01001011001011: color_data = 12'b110011110111;
		14'b01001011001100: color_data = 12'b110011110111;
		14'b01001100000000: color_data = 12'b110011110111;
		14'b01001100000001: color_data = 12'b110011110111;
		14'b01001100000010: color_data = 12'b110011110111;
		14'b01001100000011: color_data = 12'b110011110111;
		14'b01001100000100: color_data = 12'b110011110111;
		14'b01001100000101: color_data = 12'b110011110111;
		14'b01001100001011: color_data = 12'b110011110111;
		14'b01001100001100: color_data = 12'b110011110111;
		14'b01001100001101: color_data = 12'b110011110111;
		14'b01001100001110: color_data = 12'b110011110111;
		14'b01001100001111: color_data = 12'b110011110111;
		14'b01001100010000: color_data = 12'b110011110111;
		14'b01001100010110: color_data = 12'b110011110111;
		14'b01001100010111: color_data = 12'b110011110111;
		14'b01001100011000: color_data = 12'b110011110111;
		14'b01001100011001: color_data = 12'b110011110111;
		14'b01001100011010: color_data = 12'b110011110111;
		14'b01001100100001: color_data = 12'b110011110111;
		14'b01001100100010: color_data = 12'b110011110111;
		14'b01001100100011: color_data = 12'b110011110111;
		14'b01001100100100: color_data = 12'b110011110111;
		14'b01001100100101: color_data = 12'b110011110111;
		14'b01001100100110: color_data = 12'b110011110111;
		14'b01001100100111: color_data = 12'b110011110111;
		14'b01001100101000: color_data = 12'b110011110111;
		14'b01001100101001: color_data = 12'b110011110111;
		14'b01001100101010: color_data = 12'b110011110111;
		14'b01001100101011: color_data = 12'b110011110111;
		14'b01001100101100: color_data = 12'b110011110111;
		14'b01001100101101: color_data = 12'b110011110111;
		14'b01001100101110: color_data = 12'b110011110111;
		14'b01001100101111: color_data = 12'b110011110111;
		14'b01001100110000: color_data = 12'b110011110111;
		14'b01001100110110: color_data = 12'b110011110111;
		14'b01001100110111: color_data = 12'b110011110111;
		14'b01001100111000: color_data = 12'b110011110111;
		14'b01001100111001: color_data = 12'b110011110111;
		14'b01001100111010: color_data = 12'b110011110111;
		14'b01001100111011: color_data = 12'b110011110111;
		14'b01001101000001: color_data = 12'b110011110111;
		14'b01001101000010: color_data = 12'b110011110111;
		14'b01001101000011: color_data = 12'b110011110111;
		14'b01001101000100: color_data = 12'b110011110111;
		14'b01001101000101: color_data = 12'b110011110111;
		14'b01001101000110: color_data = 12'b110011110111;
		14'b01001101000111: color_data = 12'b110011110111;
		14'b01001101001000: color_data = 12'b110011110111;
		14'b01001101001001: color_data = 12'b110011110111;
		14'b01001101001010: color_data = 12'b110011110111;
		14'b01001101001011: color_data = 12'b110011110111;
		14'b01001101010001: color_data = 12'b110011110111;
		14'b01001101010010: color_data = 12'b110011110111;
		14'b01001101010011: color_data = 12'b110011110111;
		14'b01001101010100: color_data = 12'b110011110111;
		14'b01001101010101: color_data = 12'b110011110111;
		14'b01001101010110: color_data = 12'b110011110111;
		14'b01001101100001: color_data = 12'b110011110111;
		14'b01001101100010: color_data = 12'b110011110111;
		14'b01001101100011: color_data = 12'b110011110111;
		14'b01001101100100: color_data = 12'b110011110111;
		14'b01001101100101: color_data = 12'b110011110111;
		14'b01001101100110: color_data = 12'b110011110111;
		14'b01001101111100: color_data = 12'b110011110111;
		14'b01001101111101: color_data = 12'b110011110111;
		14'b01001101111110: color_data = 12'b110011110111;
		14'b01001101111111: color_data = 12'b110011110111;
		14'b01001110000000: color_data = 12'b110011110111;
		14'b01001110000001: color_data = 12'b110011110111;
		14'b01001110000111: color_data = 12'b110011110111;
		14'b01001110001000: color_data = 12'b110011110111;
		14'b01001110001001: color_data = 12'b110011110111;
		14'b01001110001010: color_data = 12'b110011110111;
		14'b01001110001011: color_data = 12'b110011110111;
		14'b01001110001100: color_data = 12'b110011110111;
		14'b01001110001101: color_data = 12'b110011110111;
		14'b01001110001110: color_data = 12'b110011110111;
		14'b01001110001111: color_data = 12'b110011110111;
		14'b01001110010000: color_data = 12'b110011110111;
		14'b01001110010001: color_data = 12'b110011110111;
		14'b01001110010010: color_data = 12'b110011110111;
		14'b01001110010011: color_data = 12'b110011110111;
		14'b01001110010100: color_data = 12'b110011110111;
		14'b01001110010101: color_data = 12'b110011110111;
		14'b01001110010110: color_data = 12'b110011110111;
		14'b01001110011101: color_data = 12'b110011110111;
		14'b01001110011110: color_data = 12'b110011110111;
		14'b01001110011111: color_data = 12'b110011110111;
		14'b01001110100000: color_data = 12'b110011110111;
		14'b01001110100001: color_data = 12'b110011110111;
		14'b01001110100010: color_data = 12'b110011110111;
		14'b01001110100011: color_data = 12'b110011110111;
		14'b01001110100100: color_data = 12'b110011110111;
		14'b01001110100101: color_data = 12'b110011110111;
		14'b01001110100110: color_data = 12'b110011110111;
		14'b01001110100111: color_data = 12'b110011110111;
		14'b01001110101000: color_data = 12'b110011110111;
		14'b01001110101001: color_data = 12'b110011110111;
		14'b01001110101010: color_data = 12'b110011110111;
		14'b01001110101011: color_data = 12'b110011110111;
		14'b01001110101100: color_data = 12'b110011110111;
		14'b01001110110010: color_data = 12'b110011110111;
		14'b01001110110011: color_data = 12'b110011110111;
		14'b01001110110100: color_data = 12'b110011110111;
		14'b01001110110101: color_data = 12'b110011110111;
		14'b01001110110110: color_data = 12'b110011110111;
		14'b01001110110111: color_data = 12'b110011110111;
		14'b01001110111000: color_data = 12'b110011110111;
		14'b01001110111001: color_data = 12'b110011110111;
		14'b01001110111010: color_data = 12'b110011110111;
		14'b01001110111011: color_data = 12'b110011110111;
		14'b01001110111100: color_data = 12'b110011110111;
		14'b01001111001000: color_data = 12'b110011110111;
		14'b01001111001001: color_data = 12'b110011110111;
		14'b01001111001010: color_data = 12'b110011110111;
		14'b01001111001011: color_data = 12'b110011110111;
		14'b01001111001100: color_data = 12'b110011110111;
		14'b01010000000000: color_data = 12'b110011110111;
		14'b01010000000001: color_data = 12'b110011110111;
		14'b01010000000010: color_data = 12'b110011110111;
		14'b01010000000011: color_data = 12'b110011110111;
		14'b01010000000100: color_data = 12'b110011110111;
		14'b01010000000101: color_data = 12'b110011110111;
		14'b01010000001011: color_data = 12'b110011110111;
		14'b01010000001100: color_data = 12'b110011110111;
		14'b01010000001101: color_data = 12'b110011110111;
		14'b01010000001110: color_data = 12'b110011110111;
		14'b01010000001111: color_data = 12'b110011110111;
		14'b01010000010000: color_data = 12'b110011110111;
		14'b01010000010110: color_data = 12'b110011110111;
		14'b01010000010111: color_data = 12'b110011110111;
		14'b01010000011000: color_data = 12'b110011110111;
		14'b01010000011001: color_data = 12'b110011110111;
		14'b01010000011010: color_data = 12'b110011110111;
		14'b01010000100001: color_data = 12'b110011110111;
		14'b01010000100010: color_data = 12'b110011110111;
		14'b01010000100011: color_data = 12'b110011110111;
		14'b01010000100100: color_data = 12'b110011110111;
		14'b01010000100101: color_data = 12'b110011110111;
		14'b01010000100110: color_data = 12'b110011110111;
		14'b01010000100111: color_data = 12'b110011110111;
		14'b01010000101000: color_data = 12'b110011110111;
		14'b01010000101001: color_data = 12'b110011110111;
		14'b01010000101010: color_data = 12'b110011110111;
		14'b01010000101011: color_data = 12'b110011110111;
		14'b01010000101100: color_data = 12'b110011110111;
		14'b01010000101101: color_data = 12'b110011110111;
		14'b01010000101110: color_data = 12'b110011110111;
		14'b01010000101111: color_data = 12'b110011110111;
		14'b01010000110000: color_data = 12'b110011110111;
		14'b01010000110110: color_data = 12'b110011110111;
		14'b01010000110111: color_data = 12'b110011110111;
		14'b01010000111000: color_data = 12'b110011110111;
		14'b01010000111001: color_data = 12'b110011110111;
		14'b01010000111010: color_data = 12'b110011110111;
		14'b01010000111011: color_data = 12'b110011110111;
		14'b01010001000001: color_data = 12'b110011110111;
		14'b01010001000010: color_data = 12'b110011110111;
		14'b01010001000011: color_data = 12'b110011110111;
		14'b01010001000100: color_data = 12'b110011110111;
		14'b01010001000101: color_data = 12'b110011110111;
		14'b01010001000110: color_data = 12'b110011110111;
		14'b01010001000111: color_data = 12'b110011110111;
		14'b01010001001000: color_data = 12'b110011110111;
		14'b01010001001001: color_data = 12'b110011110111;
		14'b01010001001010: color_data = 12'b110011110111;
		14'b01010001001011: color_data = 12'b110011110111;
		14'b01010001010001: color_data = 12'b110011110111;
		14'b01010001010010: color_data = 12'b110011110111;
		14'b01010001010011: color_data = 12'b110011110111;
		14'b01010001010100: color_data = 12'b110011110111;
		14'b01010001010101: color_data = 12'b110011110111;
		14'b01010001010110: color_data = 12'b110011110111;
		14'b01010001100001: color_data = 12'b110011110111;
		14'b01010001100010: color_data = 12'b110011110111;
		14'b01010001100011: color_data = 12'b110011110111;
		14'b01010001100100: color_data = 12'b110011110111;
		14'b01010001100101: color_data = 12'b110011110111;
		14'b01010001100110: color_data = 12'b110011110111;
		14'b01010001111100: color_data = 12'b110011110111;
		14'b01010001111101: color_data = 12'b110011110111;
		14'b01010001111110: color_data = 12'b110011110111;
		14'b01010001111111: color_data = 12'b110011110111;
		14'b01010010000000: color_data = 12'b110011110111;
		14'b01010010000001: color_data = 12'b110011110111;
		14'b01010010000111: color_data = 12'b110011110111;
		14'b01010010001000: color_data = 12'b110011110111;
		14'b01010010001001: color_data = 12'b110011110111;
		14'b01010010001010: color_data = 12'b110011110111;
		14'b01010010001011: color_data = 12'b110011110111;
		14'b01010010001100: color_data = 12'b110011110111;
		14'b01010010001101: color_data = 12'b110011110111;
		14'b01010010001110: color_data = 12'b110011110111;
		14'b01010010001111: color_data = 12'b110011110111;
		14'b01010010010000: color_data = 12'b110011110111;
		14'b01010010010001: color_data = 12'b110011110111;
		14'b01010010010010: color_data = 12'b110011110111;
		14'b01010010010011: color_data = 12'b110011110111;
		14'b01010010010100: color_data = 12'b110011110111;
		14'b01010010010101: color_data = 12'b110011110111;
		14'b01010010010110: color_data = 12'b110011110111;
		14'b01010010011101: color_data = 12'b110011110111;
		14'b01010010011110: color_data = 12'b110011110111;
		14'b01010010011111: color_data = 12'b110011110111;
		14'b01010010100000: color_data = 12'b110011110111;
		14'b01010010100001: color_data = 12'b110011110111;
		14'b01010010100010: color_data = 12'b110011110111;
		14'b01010010100011: color_data = 12'b110011110111;
		14'b01010010100100: color_data = 12'b110011110111;
		14'b01010010100101: color_data = 12'b110011110111;
		14'b01010010100110: color_data = 12'b110011110111;
		14'b01010010100111: color_data = 12'b110011110111;
		14'b01010010101000: color_data = 12'b110011110111;
		14'b01010010101001: color_data = 12'b110011110111;
		14'b01010010101010: color_data = 12'b110011110111;
		14'b01010010101011: color_data = 12'b110011110111;
		14'b01010010101100: color_data = 12'b110011110111;
		14'b01010010110010: color_data = 12'b110011110111;
		14'b01010010110011: color_data = 12'b110011110111;
		14'b01010010110100: color_data = 12'b110011110111;
		14'b01010010110101: color_data = 12'b110011110111;
		14'b01010010110110: color_data = 12'b110011110111;
		14'b01010010110111: color_data = 12'b110011110111;
		14'b01010010111000: color_data = 12'b110011110111;
		14'b01010010111001: color_data = 12'b110011110111;
		14'b01010010111010: color_data = 12'b110011110111;
		14'b01010010111011: color_data = 12'b110011110111;
		14'b01010010111100: color_data = 12'b110011110111;
		14'b01010011001000: color_data = 12'b110011110111;
		14'b01010011001001: color_data = 12'b110011110111;
		14'b01010011001010: color_data = 12'b110011110111;
		14'b01010011001011: color_data = 12'b110011110111;
		14'b01010011001100: color_data = 12'b110011110111;
		14'b01010100000000: color_data = 12'b110011110111;
		14'b01010100000001: color_data = 12'b110011110111;
		14'b01010100000010: color_data = 12'b110011110111;
		14'b01010100000011: color_data = 12'b110011110111;
		14'b01010100000100: color_data = 12'b110011110111;
		14'b01010100000101: color_data = 12'b110011110111;
		14'b01010100001011: color_data = 12'b110011110111;
		14'b01010100001100: color_data = 12'b110011110111;
		14'b01010100001101: color_data = 12'b110011110111;
		14'b01010100001110: color_data = 12'b110011110111;
		14'b01010100001111: color_data = 12'b110011110111;
		14'b01010100010000: color_data = 12'b110011110111;
		14'b01010100010110: color_data = 12'b110011110111;
		14'b01010100010111: color_data = 12'b110011110111;
		14'b01010100011000: color_data = 12'b110011110111;
		14'b01010100011001: color_data = 12'b110011110111;
		14'b01010100011010: color_data = 12'b110011110111;
		14'b01010100100001: color_data = 12'b110011110111;
		14'b01010100100010: color_data = 12'b110011110111;
		14'b01010100100011: color_data = 12'b110011110111;
		14'b01010100100100: color_data = 12'b110011110111;
		14'b01010100100101: color_data = 12'b110011110111;
		14'b01010100100110: color_data = 12'b110011110111;
		14'b01010100100111: color_data = 12'b110011110111;
		14'b01010100101000: color_data = 12'b110011110111;
		14'b01010100101001: color_data = 12'b110011110111;
		14'b01010100101010: color_data = 12'b110011110111;
		14'b01010100101011: color_data = 12'b110011110111;
		14'b01010100101100: color_data = 12'b110011110111;
		14'b01010100101101: color_data = 12'b110011110111;
		14'b01010100101110: color_data = 12'b110011110111;
		14'b01010100101111: color_data = 12'b110011110111;
		14'b01010100110000: color_data = 12'b110011110111;
		14'b01010100110110: color_data = 12'b110011110111;
		14'b01010100110111: color_data = 12'b110011110111;
		14'b01010100111000: color_data = 12'b110011110111;
		14'b01010100111001: color_data = 12'b110011110111;
		14'b01010100111010: color_data = 12'b110011110111;
		14'b01010100111011: color_data = 12'b110011110111;
		14'b01010101000001: color_data = 12'b110011110111;
		14'b01010101000010: color_data = 12'b110011110111;
		14'b01010101000011: color_data = 12'b110011110111;
		14'b01010101000100: color_data = 12'b110011110111;
		14'b01010101000101: color_data = 12'b110011110111;
		14'b01010101000110: color_data = 12'b110011110111;
		14'b01010101000111: color_data = 12'b110011110111;
		14'b01010101001000: color_data = 12'b110011110111;
		14'b01010101001001: color_data = 12'b110011110111;
		14'b01010101001010: color_data = 12'b110011110111;
		14'b01010101001011: color_data = 12'b110011110111;
		14'b01010101010001: color_data = 12'b110011110111;
		14'b01010101010010: color_data = 12'b110011110111;
		14'b01010101010011: color_data = 12'b110011110111;
		14'b01010101010100: color_data = 12'b110011110111;
		14'b01010101010101: color_data = 12'b110011110111;
		14'b01010101010110: color_data = 12'b110011110111;
		14'b01010101100001: color_data = 12'b110011110111;
		14'b01010101100010: color_data = 12'b110011110111;
		14'b01010101100011: color_data = 12'b110011110111;
		14'b01010101100100: color_data = 12'b110011110111;
		14'b01010101100101: color_data = 12'b110011110111;
		14'b01010101100110: color_data = 12'b110011110111;
		14'b01010101111100: color_data = 12'b110011110111;
		14'b01010101111101: color_data = 12'b110011110111;
		14'b01010101111110: color_data = 12'b110011110111;
		14'b01010101111111: color_data = 12'b110011110111;
		14'b01010110000000: color_data = 12'b110011110111;
		14'b01010110000001: color_data = 12'b110011110111;
		14'b01010110000111: color_data = 12'b110011110111;
		14'b01010110001000: color_data = 12'b110011110111;
		14'b01010110001001: color_data = 12'b110011110111;
		14'b01010110001010: color_data = 12'b110011110111;
		14'b01010110001011: color_data = 12'b110011110111;
		14'b01010110001100: color_data = 12'b110011110111;
		14'b01010110001101: color_data = 12'b110011110111;
		14'b01010110001110: color_data = 12'b110011110111;
		14'b01010110001111: color_data = 12'b110011110111;
		14'b01010110010000: color_data = 12'b110011110111;
		14'b01010110010001: color_data = 12'b110011110111;
		14'b01010110010010: color_data = 12'b110011110111;
		14'b01010110010011: color_data = 12'b110011110111;
		14'b01010110010100: color_data = 12'b110011110111;
		14'b01010110010101: color_data = 12'b110011110111;
		14'b01010110010110: color_data = 12'b110011110111;
		14'b01010110011101: color_data = 12'b110011110111;
		14'b01010110011110: color_data = 12'b110011110111;
		14'b01010110011111: color_data = 12'b110011110111;
		14'b01010110100000: color_data = 12'b110011110111;
		14'b01010110100001: color_data = 12'b110011110111;
		14'b01010110100010: color_data = 12'b110011110111;
		14'b01010110100011: color_data = 12'b110011110111;
		14'b01010110100100: color_data = 12'b110011110111;
		14'b01010110100101: color_data = 12'b110011110111;
		14'b01010110100110: color_data = 12'b110011110111;
		14'b01010110100111: color_data = 12'b110011110111;
		14'b01010110101000: color_data = 12'b110011110111;
		14'b01010110101001: color_data = 12'b110011110111;
		14'b01010110101010: color_data = 12'b110011110111;
		14'b01010110101011: color_data = 12'b110011110111;
		14'b01010110101100: color_data = 12'b110011110111;
		14'b01010110110010: color_data = 12'b110011110111;
		14'b01010110110011: color_data = 12'b110011110111;
		14'b01010110110100: color_data = 12'b110011110111;
		14'b01010110110101: color_data = 12'b110011110111;
		14'b01010110110110: color_data = 12'b110011110111;
		14'b01010110110111: color_data = 12'b110011110111;
		14'b01010110111000: color_data = 12'b110011110111;
		14'b01010110111001: color_data = 12'b110011110111;
		14'b01010110111010: color_data = 12'b110011110111;
		14'b01010110111011: color_data = 12'b110011110111;
		14'b01010110111100: color_data = 12'b110011110111;
		14'b01010111001000: color_data = 12'b110011110111;
		14'b01010111001001: color_data = 12'b110011110111;
		14'b01010111001010: color_data = 12'b110011110111;
		14'b01010111001011: color_data = 12'b110011110111;
		14'b01010111001100: color_data = 12'b110011110111;
		14'b01011000000000: color_data = 12'b110011110111;
		14'b01011000000001: color_data = 12'b110011110111;
		14'b01011000000010: color_data = 12'b110011110111;
		14'b01011000000011: color_data = 12'b110011110111;
		14'b01011000000100: color_data = 12'b110011110111;
		14'b01011000000101: color_data = 12'b110011110111;
		14'b01011000001011: color_data = 12'b110011110111;
		14'b01011000001100: color_data = 12'b110011110111;
		14'b01011000001101: color_data = 12'b110011110111;
		14'b01011000001110: color_data = 12'b110011110111;
		14'b01011000001111: color_data = 12'b110011110111;
		14'b01011000010000: color_data = 12'b110011110111;
		14'b01011000010110: color_data = 12'b110011110111;
		14'b01011000010111: color_data = 12'b110011110111;
		14'b01011000011000: color_data = 12'b110011110111;
		14'b01011000011001: color_data = 12'b110011110111;
		14'b01011000011010: color_data = 12'b110011110111;
		14'b01011000100001: color_data = 12'b110011110111;
		14'b01011000100010: color_data = 12'b110011110111;
		14'b01011000100011: color_data = 12'b110011110111;
		14'b01011000100100: color_data = 12'b110011110111;
		14'b01011000100101: color_data = 12'b110011110111;
		14'b01011000100110: color_data = 12'b110011110111;
		14'b01011000100111: color_data = 12'b110011110111;
		14'b01011000101000: color_data = 12'b110011110111;
		14'b01011000101001: color_data = 12'b110011110111;
		14'b01011000101010: color_data = 12'b110011110111;
		14'b01011000101011: color_data = 12'b110011110111;
		14'b01011000101100: color_data = 12'b110011110111;
		14'b01011000101101: color_data = 12'b110011110111;
		14'b01011000101110: color_data = 12'b110011110111;
		14'b01011000101111: color_data = 12'b110011110111;
		14'b01011000110000: color_data = 12'b110011110111;
		14'b01011000110110: color_data = 12'b110011110111;
		14'b01011000110111: color_data = 12'b110011110111;
		14'b01011000111000: color_data = 12'b110011110111;
		14'b01011000111001: color_data = 12'b110011110111;
		14'b01011000111010: color_data = 12'b110011110111;
		14'b01011000111011: color_data = 12'b110011110111;
		14'b01011001000001: color_data = 12'b110011110111;
		14'b01011001000010: color_data = 12'b110011110111;
		14'b01011001000011: color_data = 12'b110011110111;
		14'b01011001000100: color_data = 12'b110011110111;
		14'b01011001000101: color_data = 12'b110011110111;
		14'b01011001000110: color_data = 12'b110011110111;
		14'b01011001000111: color_data = 12'b110011110111;
		14'b01011001001000: color_data = 12'b110011110111;
		14'b01011001001001: color_data = 12'b110011110111;
		14'b01011001001010: color_data = 12'b110011110111;
		14'b01011001001011: color_data = 12'b110011110111;
		14'b01011001010001: color_data = 12'b110011110111;
		14'b01011001010010: color_data = 12'b110011110111;
		14'b01011001010011: color_data = 12'b110011110111;
		14'b01011001010100: color_data = 12'b110011110111;
		14'b01011001010101: color_data = 12'b110011110111;
		14'b01011001010110: color_data = 12'b110011110111;
		14'b01011001100001: color_data = 12'b110011110111;
		14'b01011001100010: color_data = 12'b110011110111;
		14'b01011001100011: color_data = 12'b110011110111;
		14'b01011001100100: color_data = 12'b110011110111;
		14'b01011001100101: color_data = 12'b110011110111;
		14'b01011001100110: color_data = 12'b110011110111;
		14'b01011001111100: color_data = 12'b110011110111;
		14'b01011001111101: color_data = 12'b110011110111;
		14'b01011001111110: color_data = 12'b110011110111;
		14'b01011001111111: color_data = 12'b110011110111;
		14'b01011010000000: color_data = 12'b110011110111;
		14'b01011010000001: color_data = 12'b110011110111;
		14'b01011010000111: color_data = 12'b110011110111;
		14'b01011010001000: color_data = 12'b110011110111;
		14'b01011010001001: color_data = 12'b110011110111;
		14'b01011010001010: color_data = 12'b110011110111;
		14'b01011010001011: color_data = 12'b110011110111;
		14'b01011010001100: color_data = 12'b110011110111;
		14'b01011010001101: color_data = 12'b110011110111;
		14'b01011010001110: color_data = 12'b110011110111;
		14'b01011010001111: color_data = 12'b110011110111;
		14'b01011010010000: color_data = 12'b110011110111;
		14'b01011010010001: color_data = 12'b110011110111;
		14'b01011010010010: color_data = 12'b110011110111;
		14'b01011010010011: color_data = 12'b110011110111;
		14'b01011010010100: color_data = 12'b110011110111;
		14'b01011010010101: color_data = 12'b110011110111;
		14'b01011010010110: color_data = 12'b110011110111;
		14'b01011010011101: color_data = 12'b110011110111;
		14'b01011010011110: color_data = 12'b110011110111;
		14'b01011010011111: color_data = 12'b110011110111;
		14'b01011010100000: color_data = 12'b110011110111;
		14'b01011010100001: color_data = 12'b110011110111;
		14'b01011010100010: color_data = 12'b110011110111;
		14'b01011010100011: color_data = 12'b110011110111;
		14'b01011010100100: color_data = 12'b110011110111;
		14'b01011010100101: color_data = 12'b110011110111;
		14'b01011010100110: color_data = 12'b110011110111;
		14'b01011010100111: color_data = 12'b110011110111;
		14'b01011010101000: color_data = 12'b110011110111;
		14'b01011010101001: color_data = 12'b110011110111;
		14'b01011010101010: color_data = 12'b110011110111;
		14'b01011010101011: color_data = 12'b110011110111;
		14'b01011010101100: color_data = 12'b110011110111;
		14'b01011010110010: color_data = 12'b110011110111;
		14'b01011010110011: color_data = 12'b110011110111;
		14'b01011010110100: color_data = 12'b110011110111;
		14'b01011010110101: color_data = 12'b110011110111;
		14'b01011010110110: color_data = 12'b110011110111;
		14'b01011010110111: color_data = 12'b110011110111;
		14'b01011010111000: color_data = 12'b110011110111;
		14'b01011010111001: color_data = 12'b110011110111;
		14'b01011010111010: color_data = 12'b110011110111;
		14'b01011010111011: color_data = 12'b110011110111;
		14'b01011010111100: color_data = 12'b110011110111;
		14'b01011011001000: color_data = 12'b110011110111;
		14'b01011011001001: color_data = 12'b110011110111;
		14'b01011011001010: color_data = 12'b110011110111;
		14'b01011011001011: color_data = 12'b110011110111;
		14'b01011011001100: color_data = 12'b110011110111;
		14'b01011110100111: color_data = 12'b110011110111;
		14'b01011110101000: color_data = 12'b110011110111;
		14'b01011110101001: color_data = 12'b110011110111;
		14'b01011110101010: color_data = 12'b110011110111;
		14'b01011110101011: color_data = 12'b110011110111;
		14'b01011110101100: color_data = 12'b110011110111;
		14'b01100010100111: color_data = 12'b110011110111;
		14'b01100010101000: color_data = 12'b110011110111;
		14'b01100010101001: color_data = 12'b110011110111;
		14'b01100010101010: color_data = 12'b110011110111;
		14'b01100010101011: color_data = 12'b110011110111;
		14'b01100010101100: color_data = 12'b110011110111;
		14'b01100110100111: color_data = 12'b110011110111;
		14'b01100110101000: color_data = 12'b110011110111;
		14'b01100110101001: color_data = 12'b110011110111;
		14'b01100110101010: color_data = 12'b110011110111;
		14'b01100110101011: color_data = 12'b110011110111;
		14'b01100110101100: color_data = 12'b110011110111;
		14'b01101010100111: color_data = 12'b110011110111;
		14'b01101010101000: color_data = 12'b110011110111;
		14'b01101010101001: color_data = 12'b110011110111;
		14'b01101010101010: color_data = 12'b110011110111;
		14'b01101010101011: color_data = 12'b110011110111;
		14'b01101010101100: color_data = 12'b110011110111;
		14'b01101110100111: color_data = 12'b110011110111;
		14'b01101110101000: color_data = 12'b110011110111;
		14'b01101110101001: color_data = 12'b110011110111;
		14'b01101110101010: color_data = 12'b110011110111;
		14'b01101110101011: color_data = 12'b110011110111;
		14'b01101110101100: color_data = 12'b110011110111;
		14'b01110010011101: color_data = 12'b110011110111;
		14'b01110010011110: color_data = 12'b110011110111;
		14'b01110010011111: color_data = 12'b110011110111;
		14'b01110010100000: color_data = 12'b110011110111;
		14'b01110010100001: color_data = 12'b110011110111;
		14'b01110010100010: color_data = 12'b110011110111;
		14'b01110010100011: color_data = 12'b110011110111;
		14'b01110010100100: color_data = 12'b110011110111;
		14'b01110010100101: color_data = 12'b110011110111;
		14'b01110010100110: color_data = 12'b110011110111;
		14'b01110010100111: color_data = 12'b110011110111;
		14'b01110010101000: color_data = 12'b110011110111;
		14'b01110010101001: color_data = 12'b110011110111;
		14'b01110010101010: color_data = 12'b110011110111;
		14'b01110010101011: color_data = 12'b110011110111;
		14'b01110010101100: color_data = 12'b110011110111;
		14'b01110110011101: color_data = 12'b110011110111;
		14'b01110110011110: color_data = 12'b110011110111;
		14'b01110110011111: color_data = 12'b110011110111;
		14'b01110110100000: color_data = 12'b110011110111;
		14'b01110110100001: color_data = 12'b110011110111;
		14'b01110110100010: color_data = 12'b110011110111;
		14'b01110110100011: color_data = 12'b110011110111;
		14'b01110110100100: color_data = 12'b110011110111;
		14'b01110110100101: color_data = 12'b110011110111;
		14'b01110110100110: color_data = 12'b110011110111;
		14'b01110110100111: color_data = 12'b110011110111;
		14'b01110110101000: color_data = 12'b110011110111;
		14'b01110110101001: color_data = 12'b110011110111;
		14'b01110110101010: color_data = 12'b110011110111;
		14'b01110110101011: color_data = 12'b110011110111;
		14'b01110110101100: color_data = 12'b110011110111;
		14'b01111010011101: color_data = 12'b110011110111;
		14'b01111010011110: color_data = 12'b110011110111;
		14'b01111010011111: color_data = 12'b110011110111;
		14'b01111010100000: color_data = 12'b110011110111;
		14'b01111010100001: color_data = 12'b110011110111;
		14'b01111010100010: color_data = 12'b110011110111;
		14'b01111010100011: color_data = 12'b110011110111;
		14'b01111010100100: color_data = 12'b110011110111;
		14'b01111010100101: color_data = 12'b110011110111;
		14'b01111010100110: color_data = 12'b110011110111;
		14'b01111010100111: color_data = 12'b110011110111;
		14'b01111010101000: color_data = 12'b110011110111;
		14'b01111010101001: color_data = 12'b110011110111;
		14'b01111010101010: color_data = 12'b110011110111;
		14'b01111010101011: color_data = 12'b110011110111;
		14'b01111010101100: color_data = 12'b110011110111;
		14'b01111110011101: color_data = 12'b110011110111;
		14'b01111110011110: color_data = 12'b110011110111;
		14'b01111110011111: color_data = 12'b110011110111;
		14'b01111110100000: color_data = 12'b110011110111;
		14'b01111110100001: color_data = 12'b110011110111;
		14'b01111110100010: color_data = 12'b110011110111;
		14'b01111110100011: color_data = 12'b110011110111;
		14'b01111110100100: color_data = 12'b110011110111;
		14'b01111110100101: color_data = 12'b110011110111;
		14'b01111110100110: color_data = 12'b110011110111;
		14'b01111110100111: color_data = 12'b110011110111;
		14'b01111110101000: color_data = 12'b110011110111;
		14'b01111110101001: color_data = 12'b110011110111;
		14'b01111110101010: color_data = 12'b110011110111;
		14'b01111110101011: color_data = 12'b110011110111;
		14'b01111110101100: color_data = 12'b110011110111;
		14'b10000010011101: color_data = 12'b110011110111;
		14'b10000010011110: color_data = 12'b110011110111;
		14'b10000010011111: color_data = 12'b110011110111;
		14'b10000010100000: color_data = 12'b110011110111;
		14'b10000010100001: color_data = 12'b110011110111;
		14'b10000010100010: color_data = 12'b110011110111;
		14'b10000010100011: color_data = 12'b110011110111;
		14'b10000010100100: color_data = 12'b110011110111;
		14'b10000010100101: color_data = 12'b110011110111;
		14'b10000010100110: color_data = 12'b110011110111;
		14'b10000010100111: color_data = 12'b110011110111;
		14'b10000010101000: color_data = 12'b110011110111;
		14'b10000010101001: color_data = 12'b110011110111;
		14'b10000010101010: color_data = 12'b110011110111;
		14'b10000010101011: color_data = 12'b110011110111;
		14'b10000010101100: color_data = 12'b110011110111;

		default:color_data = 12'd0;
	endcase
endmodule
