`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.01.2025 16:24:33
// Design Name: 
// Module Name: single_text_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module single_text_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [7:0] col,
		output reg [11:0] color_data
	);

	
    (* rom_style = "block" *)
	//signal declaration
	reg [5:0] row_reg;
	reg [7:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		14'b00000000000000: color_data = 12'b110011110111;
		14'b00000000000001: color_data = 12'b110011110111;
		14'b00000000000010: color_data = 12'b110011110111;
		14'b00000000000011: color_data = 12'b110011110111;
		14'b00000000000100: color_data = 12'b110011110111;
		14'b00000000000101: color_data = 12'b110011110111;
		14'b00000000000110: color_data = 12'b110011110111;
		14'b00000000000111: color_data = 12'b110011110111;
		14'b00000000001000: color_data = 12'b110011110111;
		14'b00000000001001: color_data = 12'b110011110111;
		14'b00000000001010: color_data = 12'b110011110111;
		14'b00000000001011: color_data = 12'b110011110111;
		14'b00000000001100: color_data = 12'b110011110111;
		14'b00000000001101: color_data = 12'b110011110111;
		14'b00000000001110: color_data = 12'b110011110111;
		14'b00000000001111: color_data = 12'b110011110111;
		14'b00000000010000: color_data = 12'b110011110111;
		14'b00000000010001: color_data = 12'b110011110111;
		14'b00000000010010: color_data = 12'b110011110111;
		14'b00000000010011: color_data = 12'b110011110111;
		14'b00000000011001: color_data = 12'b110011110111;
		14'b00000000011010: color_data = 12'b110011110111;
		14'b00000000011011: color_data = 12'b110011110111;
		14'b00000000011100: color_data = 12'b110011110111;
		14'b00000000011101: color_data = 12'b110011110111;
		14'b00000001001010: color_data = 12'b110011110111;
		14'b00000001001011: color_data = 12'b110011110111;
		14'b00000001001100: color_data = 12'b110011110111;
		14'b00000001001101: color_data = 12'b110011110111;
		14'b00000001001110: color_data = 12'b110011110111;
		14'b00000001101100: color_data = 12'b110011110111;
		14'b00000001101101: color_data = 12'b110011110111;
		14'b00000001101110: color_data = 12'b110011110111;
		14'b00000001101111: color_data = 12'b110011110111;
		14'b00000001110000: color_data = 12'b110011110111;
		14'b00000001110001: color_data = 12'b110011110111;
		14'b00000001110010: color_data = 12'b110011110111;
		14'b00000001110011: color_data = 12'b110011110111;
		14'b00000001110100: color_data = 12'b110011110111;
		14'b00000001110101: color_data = 12'b110011110111;
		14'b00000001110110: color_data = 12'b110011110111;
		14'b00000001110111: color_data = 12'b110011110111;
		14'b00000001111000: color_data = 12'b110011110111;
		14'b00000001111001: color_data = 12'b110011110111;
		14'b00000001111010: color_data = 12'b110011110111;
		14'b00000001111011: color_data = 12'b110011110111;
		14'b00000001111100: color_data = 12'b110011110111;
		14'b00000001111101: color_data = 12'b110011110111;
		14'b00000001111110: color_data = 12'b110011110111;
		14'b00000010000100: color_data = 12'b110011110111;
		14'b00000010000101: color_data = 12'b110011110111;
		14'b00000010000110: color_data = 12'b110011110111;
		14'b00000010000111: color_data = 12'b110011110111;
		14'b00000010001000: color_data = 12'b110011110111;
		14'b00000100000000: color_data = 12'b110011110111;
		14'b00000100000001: color_data = 12'b110011110111;
		14'b00000100000010: color_data = 12'b110011110111;
		14'b00000100000011: color_data = 12'b110011110111;
		14'b00000100000100: color_data = 12'b110011110111;
		14'b00000100000101: color_data = 12'b110011110111;
		14'b00000100000110: color_data = 12'b110011110111;
		14'b00000100000111: color_data = 12'b110011110111;
		14'b00000100001000: color_data = 12'b110011110111;
		14'b00000100001001: color_data = 12'b110011110111;
		14'b00000100001010: color_data = 12'b110011110111;
		14'b00000100001011: color_data = 12'b110011110111;
		14'b00000100001100: color_data = 12'b110011110111;
		14'b00000100001101: color_data = 12'b110011110111;
		14'b00000100001110: color_data = 12'b110011110111;
		14'b00000100001111: color_data = 12'b110011110111;
		14'b00000100010000: color_data = 12'b110011110111;
		14'b00000100010001: color_data = 12'b110011110111;
		14'b00000100010010: color_data = 12'b110011110111;
		14'b00000100010011: color_data = 12'b110011110111;
		14'b00000100011001: color_data = 12'b110011110111;
		14'b00000100011010: color_data = 12'b110011110111;
		14'b00000100011011: color_data = 12'b110011110111;
		14'b00000100011100: color_data = 12'b110011110111;
		14'b00000100011101: color_data = 12'b110011110111;
		14'b00000101001010: color_data = 12'b110011110111;
		14'b00000101001011: color_data = 12'b110011110111;
		14'b00000101001100: color_data = 12'b110011110111;
		14'b00000101001101: color_data = 12'b110011110111;
		14'b00000101001110: color_data = 12'b110011110111;
		14'b00000101101100: color_data = 12'b110011110111;
		14'b00000101101101: color_data = 12'b110011110111;
		14'b00000101101110: color_data = 12'b110011110111;
		14'b00000101101111: color_data = 12'b110011110111;
		14'b00000101110000: color_data = 12'b110011110111;
		14'b00000101110001: color_data = 12'b110011110111;
		14'b00000101110010: color_data = 12'b110011110111;
		14'b00000101110011: color_data = 12'b110011110111;
		14'b00000101110100: color_data = 12'b110011110111;
		14'b00000101110101: color_data = 12'b110011110111;
		14'b00000101110110: color_data = 12'b110011110111;
		14'b00000101110111: color_data = 12'b110011110111;
		14'b00000101111000: color_data = 12'b110011110111;
		14'b00000101111001: color_data = 12'b110011110111;
		14'b00000101111010: color_data = 12'b110011110111;
		14'b00000101111011: color_data = 12'b110011110111;
		14'b00000101111100: color_data = 12'b110011110111;
		14'b00000101111101: color_data = 12'b110011110111;
		14'b00000101111110: color_data = 12'b110011110111;
		14'b00000110000100: color_data = 12'b110011110111;
		14'b00000110000101: color_data = 12'b110011110111;
		14'b00000110000110: color_data = 12'b110011110111;
		14'b00000110000111: color_data = 12'b110011110111;
		14'b00000110001000: color_data = 12'b110011110111;
		14'b00001000000000: color_data = 12'b110011110111;
		14'b00001000000001: color_data = 12'b110011110111;
		14'b00001000000010: color_data = 12'b110011110111;
		14'b00001000000011: color_data = 12'b110011110111;
		14'b00001000000100: color_data = 12'b110011110111;
		14'b00001000000101: color_data = 12'b110011110111;
		14'b00001000000110: color_data = 12'b110011110111;
		14'b00001000000111: color_data = 12'b110011110111;
		14'b00001000001000: color_data = 12'b110011110111;
		14'b00001000001001: color_data = 12'b110011110111;
		14'b00001000001010: color_data = 12'b110011110111;
		14'b00001000001011: color_data = 12'b110011110111;
		14'b00001000001100: color_data = 12'b110011110111;
		14'b00001000001101: color_data = 12'b110011110111;
		14'b00001000001110: color_data = 12'b110011110111;
		14'b00001000001111: color_data = 12'b110011110111;
		14'b00001000010000: color_data = 12'b110011110111;
		14'b00001000010001: color_data = 12'b110011110111;
		14'b00001000010010: color_data = 12'b110011110111;
		14'b00001000010011: color_data = 12'b110011110111;
		14'b00001000011001: color_data = 12'b110011110111;
		14'b00001000011010: color_data = 12'b110011110111;
		14'b00001000011011: color_data = 12'b110011110111;
		14'b00001000011100: color_data = 12'b110011110111;
		14'b00001000011101: color_data = 12'b110011110111;
		14'b00001001001010: color_data = 12'b110011110111;
		14'b00001001001011: color_data = 12'b110011110111;
		14'b00001001001100: color_data = 12'b110011110111;
		14'b00001001001101: color_data = 12'b110011110111;
		14'b00001001001110: color_data = 12'b110011110111;
		14'b00001001101100: color_data = 12'b110011110111;
		14'b00001001101101: color_data = 12'b110011110111;
		14'b00001001101110: color_data = 12'b110011110111;
		14'b00001001101111: color_data = 12'b110011110111;
		14'b00001001110000: color_data = 12'b110011110111;
		14'b00001001110001: color_data = 12'b110011110111;
		14'b00001001110010: color_data = 12'b110011110111;
		14'b00001001110011: color_data = 12'b110011110111;
		14'b00001001110100: color_data = 12'b110011110111;
		14'b00001001110101: color_data = 12'b110011110111;
		14'b00001001110110: color_data = 12'b110011110111;
		14'b00001001110111: color_data = 12'b110011110111;
		14'b00001001111000: color_data = 12'b110011110111;
		14'b00001001111001: color_data = 12'b110011110111;
		14'b00001001111010: color_data = 12'b110011110111;
		14'b00001001111011: color_data = 12'b110011110111;
		14'b00001001111100: color_data = 12'b110011110111;
		14'b00001001111101: color_data = 12'b110011110111;
		14'b00001001111110: color_data = 12'b110011110111;
		14'b00001010000100: color_data = 12'b110011110111;
		14'b00001010000101: color_data = 12'b110011110111;
		14'b00001010000110: color_data = 12'b110011110111;
		14'b00001010000111: color_data = 12'b110011110111;
		14'b00001010001000: color_data = 12'b110011110111;
		14'b00001100000000: color_data = 12'b110011110111;
		14'b00001100000001: color_data = 12'b110011110111;
		14'b00001100000010: color_data = 12'b110011110111;
		14'b00001100000011: color_data = 12'b110011110111;
		14'b00001100000100: color_data = 12'b110011110111;
		14'b00001100000101: color_data = 12'b110011110111;
		14'b00001100000110: color_data = 12'b110011110111;
		14'b00001100000111: color_data = 12'b110011110111;
		14'b00001100001000: color_data = 12'b110011110111;
		14'b00001100001001: color_data = 12'b110011110111;
		14'b00001100001010: color_data = 12'b110011110111;
		14'b00001100001011: color_data = 12'b110011110111;
		14'b00001100001100: color_data = 12'b110011110111;
		14'b00001100001101: color_data = 12'b110011110111;
		14'b00001100001110: color_data = 12'b110011110111;
		14'b00001100001111: color_data = 12'b110011110111;
		14'b00001100010000: color_data = 12'b110011110111;
		14'b00001100010001: color_data = 12'b110011110111;
		14'b00001100010010: color_data = 12'b110011110111;
		14'b00001100010011: color_data = 12'b110011110111;
		14'b00001100011001: color_data = 12'b110011110111;
		14'b00001100011010: color_data = 12'b110011110111;
		14'b00001100011011: color_data = 12'b110011110111;
		14'b00001100011100: color_data = 12'b110011110111;
		14'b00001100011101: color_data = 12'b110011110111;
		14'b00001101001010: color_data = 12'b110011110111;
		14'b00001101001011: color_data = 12'b110011110111;
		14'b00001101001100: color_data = 12'b110011110111;
		14'b00001101001101: color_data = 12'b110011110111;
		14'b00001101001110: color_data = 12'b110011110111;
		14'b00001101101100: color_data = 12'b110011110111;
		14'b00001101101101: color_data = 12'b110011110111;
		14'b00001101101110: color_data = 12'b110011110111;
		14'b00001101101111: color_data = 12'b110011110111;
		14'b00001101110000: color_data = 12'b110011110111;
		14'b00001101110001: color_data = 12'b110011110111;
		14'b00001101110010: color_data = 12'b110011110111;
		14'b00001101110011: color_data = 12'b110011110111;
		14'b00001101110100: color_data = 12'b110011110111;
		14'b00001101110101: color_data = 12'b110011110111;
		14'b00001101110110: color_data = 12'b110011110111;
		14'b00001101110111: color_data = 12'b110011110111;
		14'b00001101111000: color_data = 12'b110011110111;
		14'b00001101111001: color_data = 12'b110011110111;
		14'b00001101111010: color_data = 12'b110011110111;
		14'b00001101111011: color_data = 12'b110011110111;
		14'b00001101111100: color_data = 12'b110011110111;
		14'b00001101111101: color_data = 12'b110011110111;
		14'b00001101111110: color_data = 12'b110011110111;
		14'b00001110000100: color_data = 12'b110011110111;
		14'b00001110000101: color_data = 12'b110011110111;
		14'b00001110000110: color_data = 12'b110011110111;
		14'b00001110000111: color_data = 12'b110011110111;
		14'b00001110001000: color_data = 12'b110011110111;
		14'b00010000000000: color_data = 12'b110011110111;
		14'b00010000000001: color_data = 12'b110011110111;
		14'b00010000000010: color_data = 12'b110011110111;
		14'b00010000000011: color_data = 12'b110011110111;
		14'b00010000000100: color_data = 12'b110011110111;
		14'b00010000000101: color_data = 12'b110011110111;
		14'b00010000000110: color_data = 12'b110011110111;
		14'b00010000000111: color_data = 12'b110011110111;
		14'b00010000001000: color_data = 12'b110011110111;
		14'b00010000001001: color_data = 12'b110011110111;
		14'b00010000001010: color_data = 12'b110011110111;
		14'b00010000001011: color_data = 12'b110011110111;
		14'b00010000001100: color_data = 12'b110011110111;
		14'b00010000001101: color_data = 12'b110011110111;
		14'b00010000001110: color_data = 12'b110011110111;
		14'b00010000001111: color_data = 12'b110011110111;
		14'b00010000010000: color_data = 12'b110011110111;
		14'b00010000010001: color_data = 12'b110011110111;
		14'b00010000010010: color_data = 12'b110011110111;
		14'b00010000010011: color_data = 12'b110011110111;
		14'b00010000011001: color_data = 12'b110011110111;
		14'b00010000011010: color_data = 12'b110011110111;
		14'b00010000011011: color_data = 12'b110011110111;
		14'b00010000011100: color_data = 12'b110011110111;
		14'b00010000011101: color_data = 12'b110011110111;
		14'b00010001001010: color_data = 12'b110011110111;
		14'b00010001001011: color_data = 12'b110011110111;
		14'b00010001001100: color_data = 12'b110011110111;
		14'b00010001001101: color_data = 12'b110011110111;
		14'b00010001001110: color_data = 12'b110011110111;
		14'b00010001101100: color_data = 12'b110011110111;
		14'b00010001101101: color_data = 12'b110011110111;
		14'b00010001101110: color_data = 12'b110011110111;
		14'b00010001101111: color_data = 12'b110011110111;
		14'b00010001110000: color_data = 12'b110011110111;
		14'b00010001110001: color_data = 12'b110011110111;
		14'b00010001110010: color_data = 12'b110011110111;
		14'b00010001110011: color_data = 12'b110011110111;
		14'b00010001110100: color_data = 12'b110011110111;
		14'b00010001110101: color_data = 12'b110011110111;
		14'b00010001110110: color_data = 12'b110011110111;
		14'b00010001110111: color_data = 12'b110011110111;
		14'b00010001111000: color_data = 12'b110011110111;
		14'b00010001111001: color_data = 12'b110011110111;
		14'b00010001111010: color_data = 12'b110011110111;
		14'b00010001111011: color_data = 12'b110011110111;
		14'b00010001111100: color_data = 12'b110011110111;
		14'b00010001111101: color_data = 12'b110011110111;
		14'b00010001111110: color_data = 12'b110011110111;
		14'b00010010000100: color_data = 12'b110011110111;
		14'b00010010000101: color_data = 12'b110011110111;
		14'b00010010000110: color_data = 12'b110011110111;
		14'b00010010000111: color_data = 12'b110011110111;
		14'b00010010001000: color_data = 12'b110011110111;
		14'b00010100000000: color_data = 12'b110011110111;
		14'b00010100000001: color_data = 12'b110011110111;
		14'b00010100000010: color_data = 12'b110011110111;
		14'b00010100000011: color_data = 12'b110011110111;
		14'b00010100000100: color_data = 12'b110011110111;
		14'b00010101001010: color_data = 12'b110011110111;
		14'b00010101001011: color_data = 12'b110011110111;
		14'b00010101001100: color_data = 12'b110011110111;
		14'b00010101001101: color_data = 12'b110011110111;
		14'b00010101001110: color_data = 12'b110011110111;
		14'b00010101101100: color_data = 12'b110011110111;
		14'b00010101101101: color_data = 12'b110011110111;
		14'b00010101101110: color_data = 12'b110011110111;
		14'b00010101101111: color_data = 12'b110011110111;
		14'b00010101110000: color_data = 12'b110011110111;
		14'b00010101111011: color_data = 12'b110011110111;
		14'b00010101111100: color_data = 12'b110011110111;
		14'b00010101111101: color_data = 12'b110011110111;
		14'b00010101111110: color_data = 12'b110011110111;
		14'b00010110000100: color_data = 12'b110011110111;
		14'b00010110000101: color_data = 12'b110011110111;
		14'b00010110000110: color_data = 12'b110011110111;
		14'b00010110000111: color_data = 12'b110011110111;
		14'b00010110001000: color_data = 12'b110011110111;
		14'b00011000000000: color_data = 12'b110011110111;
		14'b00011000000001: color_data = 12'b110011110111;
		14'b00011000000010: color_data = 12'b110011110111;
		14'b00011000000011: color_data = 12'b110011110111;
		14'b00011000000100: color_data = 12'b110011110111;
		14'b00011001001010: color_data = 12'b110011110111;
		14'b00011001001011: color_data = 12'b110011110111;
		14'b00011001001100: color_data = 12'b110011110111;
		14'b00011001001101: color_data = 12'b110011110111;
		14'b00011001001110: color_data = 12'b110011110111;
		14'b00011001101100: color_data = 12'b110011110111;
		14'b00011001101101: color_data = 12'b110011110111;
		14'b00011001101110: color_data = 12'b110011110111;
		14'b00011001101111: color_data = 12'b110011110111;
		14'b00011001110000: color_data = 12'b110011110111;
		14'b00011001111011: color_data = 12'b110011110111;
		14'b00011001111100: color_data = 12'b110011110111;
		14'b00011001111101: color_data = 12'b110011110111;
		14'b00011001111110: color_data = 12'b110011110111;
		14'b00011010000100: color_data = 12'b110011110111;
		14'b00011010000101: color_data = 12'b110011110111;
		14'b00011010000110: color_data = 12'b110011110111;
		14'b00011010000111: color_data = 12'b110011110111;
		14'b00011010001000: color_data = 12'b110011110111;
		14'b00011100000000: color_data = 12'b110011110111;
		14'b00011100000001: color_data = 12'b110011110111;
		14'b00011100000010: color_data = 12'b110011110111;
		14'b00011100000011: color_data = 12'b110011110111;
		14'b00011100000100: color_data = 12'b110011110111;
		14'b00011101001010: color_data = 12'b110011110111;
		14'b00011101001011: color_data = 12'b110011110111;
		14'b00011101001100: color_data = 12'b110011110111;
		14'b00011101001101: color_data = 12'b110011110111;
		14'b00011101001110: color_data = 12'b110011110111;
		14'b00011101101100: color_data = 12'b110011110111;
		14'b00011101101101: color_data = 12'b110011110111;
		14'b00011101101110: color_data = 12'b110011110111;
		14'b00011101101111: color_data = 12'b110011110111;
		14'b00011101110000: color_data = 12'b110011110111;
		14'b00011101111011: color_data = 12'b110011110111;
		14'b00011101111100: color_data = 12'b110011110111;
		14'b00011101111101: color_data = 12'b110011110111;
		14'b00011101111110: color_data = 12'b110011110111;
		14'b00011110000100: color_data = 12'b110011110111;
		14'b00011110000101: color_data = 12'b110011110111;
		14'b00011110000110: color_data = 12'b110011110111;
		14'b00011110000111: color_data = 12'b110011110111;
		14'b00011110001000: color_data = 12'b110011110111;
		14'b00100000000000: color_data = 12'b110011110111;
		14'b00100000000001: color_data = 12'b110011110111;
		14'b00100000000010: color_data = 12'b110011110111;
		14'b00100000000011: color_data = 12'b110011110111;
		14'b00100000000100: color_data = 12'b110011110111;
		14'b00100001001010: color_data = 12'b110011110111;
		14'b00100001001011: color_data = 12'b110011110111;
		14'b00100001001100: color_data = 12'b110011110111;
		14'b00100001001101: color_data = 12'b110011110111;
		14'b00100001001110: color_data = 12'b110011110111;
		14'b00100001101100: color_data = 12'b110011110111;
		14'b00100001101101: color_data = 12'b110011110111;
		14'b00100001101110: color_data = 12'b110011110111;
		14'b00100001101111: color_data = 12'b110011110111;
		14'b00100001110000: color_data = 12'b110011110111;
		14'b00100001111011: color_data = 12'b110011110111;
		14'b00100001111100: color_data = 12'b110011110111;
		14'b00100001111101: color_data = 12'b110011110111;
		14'b00100001111110: color_data = 12'b110011110111;
		14'b00100010000100: color_data = 12'b110011110111;
		14'b00100010000101: color_data = 12'b110011110111;
		14'b00100010000110: color_data = 12'b110011110111;
		14'b00100010000111: color_data = 12'b110011110111;
		14'b00100010001000: color_data = 12'b110011110111;
		14'b00100100000000: color_data = 12'b110011110111;
		14'b00100100000001: color_data = 12'b110011110111;
		14'b00100100000010: color_data = 12'b110011110111;
		14'b00100100000011: color_data = 12'b110011110111;
		14'b00100100000100: color_data = 12'b110011110111;
		14'b00100100000101: color_data = 12'b110011110111;
		14'b00100100000110: color_data = 12'b110011110111;
		14'b00100100000111: color_data = 12'b110011110111;
		14'b00100100001000: color_data = 12'b110011110111;
		14'b00100100001001: color_data = 12'b110011110111;
		14'b00100100001010: color_data = 12'b110011110111;
		14'b00100100001011: color_data = 12'b110011110111;
		14'b00100100001100: color_data = 12'b110011110111;
		14'b00100100001101: color_data = 12'b110011110111;
		14'b00100100001110: color_data = 12'b110011110111;
		14'b00100100001111: color_data = 12'b110011110111;
		14'b00100100010000: color_data = 12'b110011110111;
		14'b00100100010001: color_data = 12'b110011110111;
		14'b00100100010010: color_data = 12'b110011110111;
		14'b00100100010011: color_data = 12'b110011110111;
		14'b00100100011001: color_data = 12'b110011110111;
		14'b00100100011010: color_data = 12'b110011110111;
		14'b00100100011011: color_data = 12'b110011110111;
		14'b00100100011100: color_data = 12'b110011110111;
		14'b00100100011101: color_data = 12'b110011110111;
		14'b00100100100011: color_data = 12'b110011110111;
		14'b00100100100100: color_data = 12'b110011110111;
		14'b00100100100101: color_data = 12'b110011110111;
		14'b00100100100110: color_data = 12'b110011110111;
		14'b00100100100111: color_data = 12'b110011110111;
		14'b00100100101000: color_data = 12'b110011110111;
		14'b00100100101001: color_data = 12'b110011110111;
		14'b00100100101010: color_data = 12'b110011110111;
		14'b00100100101011: color_data = 12'b110011110111;
		14'b00100100101100: color_data = 12'b110011110111;
		14'b00100100101101: color_data = 12'b110011110111;
		14'b00100100101110: color_data = 12'b110011110111;
		14'b00100100101111: color_data = 12'b110011110111;
		14'b00100100110000: color_data = 12'b110011110111;
		14'b00100100110110: color_data = 12'b110011110111;
		14'b00100100110111: color_data = 12'b110011110111;
		14'b00100100111000: color_data = 12'b110011110111;
		14'b00100100111001: color_data = 12'b110011110111;
		14'b00100100111010: color_data = 12'b110011110111;
		14'b00100100111011: color_data = 12'b110011110111;
		14'b00100100111100: color_data = 12'b110011110111;
		14'b00100100111101: color_data = 12'b110011110111;
		14'b00100100111110: color_data = 12'b110011110111;
		14'b00100100111111: color_data = 12'b110011110111;
		14'b00100101000000: color_data = 12'b110011110111;
		14'b00100101000001: color_data = 12'b110011110111;
		14'b00100101000010: color_data = 12'b110011110111;
		14'b00100101000011: color_data = 12'b110011110111;
		14'b00100101000100: color_data = 12'b110011110111;
		14'b00100101001010: color_data = 12'b110011110111;
		14'b00100101001011: color_data = 12'b110011110111;
		14'b00100101001100: color_data = 12'b110011110111;
		14'b00100101001101: color_data = 12'b110011110111;
		14'b00100101001110: color_data = 12'b110011110111;
		14'b00100101010100: color_data = 12'b110011110111;
		14'b00100101010101: color_data = 12'b110011110111;
		14'b00100101010110: color_data = 12'b110011110111;
		14'b00100101010111: color_data = 12'b110011110111;
		14'b00100101011000: color_data = 12'b110011110111;
		14'b00100101011001: color_data = 12'b110011110111;
		14'b00100101011010: color_data = 12'b110011110111;
		14'b00100101011011: color_data = 12'b110011110111;
		14'b00100101011100: color_data = 12'b110011110111;
		14'b00100101011101: color_data = 12'b110011110111;
		14'b00100101011110: color_data = 12'b110011110111;
		14'b00100101011111: color_data = 12'b110011110111;
		14'b00100101100000: color_data = 12'b110011110111;
		14'b00100101100001: color_data = 12'b110011110111;
		14'b00100101101100: color_data = 12'b110011110111;
		14'b00100101101101: color_data = 12'b110011110111;
		14'b00100101101110: color_data = 12'b110011110111;
		14'b00100101101111: color_data = 12'b110011110111;
		14'b00100101110000: color_data = 12'b110011110111;
		14'b00100101110001: color_data = 12'b110011110111;
		14'b00100101110010: color_data = 12'b110011110111;
		14'b00100101110011: color_data = 12'b110011110111;
		14'b00100101110100: color_data = 12'b110011110111;
		14'b00100101110101: color_data = 12'b110011110111;
		14'b00100101110110: color_data = 12'b110011110111;
		14'b00100101110111: color_data = 12'b110011110111;
		14'b00100101111000: color_data = 12'b110011110111;
		14'b00100101111001: color_data = 12'b110011110111;
		14'b00100101111010: color_data = 12'b110011110111;
		14'b00100101111011: color_data = 12'b110011110111;
		14'b00100101111100: color_data = 12'b110011110111;
		14'b00100101111101: color_data = 12'b110011110111;
		14'b00100101111110: color_data = 12'b110011110111;
		14'b00100110000100: color_data = 12'b110011110111;
		14'b00100110000101: color_data = 12'b110011110111;
		14'b00100110000110: color_data = 12'b110011110111;
		14'b00100110000111: color_data = 12'b110011110111;
		14'b00100110001000: color_data = 12'b110011110111;
		14'b00100110010011: color_data = 12'b110011110111;
		14'b00100110010100: color_data = 12'b110011110111;
		14'b00100110010101: color_data = 12'b110011110111;
		14'b00100110010110: color_data = 12'b110011110111;
		14'b00100110010111: color_data = 12'b110011110111;
		14'b00100110011000: color_data = 12'b110011110111;
		14'b00100110011001: color_data = 12'b110011110111;
		14'b00100110011010: color_data = 12'b110011110111;
		14'b00100110011011: color_data = 12'b110011110111;
		14'b00100110011100: color_data = 12'b110011110111;
		14'b00100110100010: color_data = 12'b110011110111;
		14'b00100110100011: color_data = 12'b110011110111;
		14'b00100110100100: color_data = 12'b110011110111;
		14'b00100110100101: color_data = 12'b110011110111;
		14'b00100110100110: color_data = 12'b110011110111;
		14'b00100110101011: color_data = 12'b110011110111;
		14'b00100110101100: color_data = 12'b110011110111;
		14'b00100110101101: color_data = 12'b110011110111;
		14'b00100110101110: color_data = 12'b110011110111;
		14'b00100110101111: color_data = 12'b110011110111;
		14'b00100110110101: color_data = 12'b110011110111;
		14'b00100110110110: color_data = 12'b110011110111;
		14'b00100110110111: color_data = 12'b110011110111;
		14'b00100110111000: color_data = 12'b110011110111;
		14'b00100110111001: color_data = 12'b110011110111;
		14'b00100110111010: color_data = 12'b110011110111;
		14'b00100110111011: color_data = 12'b110011110111;
		14'b00100110111100: color_data = 12'b110011110111;
		14'b00100110111101: color_data = 12'b110011110111;
		14'b00100110111110: color_data = 12'b110011110111;
		14'b00100110111111: color_data = 12'b110011110111;
		14'b00100111000000: color_data = 12'b110011110111;
		14'b00100111000001: color_data = 12'b110011110111;
		14'b00100111000010: color_data = 12'b110011110111;
		14'b00100111000011: color_data = 12'b110011110111;
		14'b00100111001001: color_data = 12'b110011110111;
		14'b00100111001010: color_data = 12'b110011110111;
		14'b00100111001011: color_data = 12'b110011110111;
		14'b00100111001100: color_data = 12'b110011110111;
		14'b00100111001101: color_data = 12'b110011110111;
		14'b00100111001110: color_data = 12'b110011110111;
		14'b00100111001111: color_data = 12'b110011110111;
		14'b00100111010000: color_data = 12'b110011110111;
		14'b00100111010001: color_data = 12'b110011110111;
		14'b00101000000000: color_data = 12'b110011110111;
		14'b00101000000001: color_data = 12'b110011110111;
		14'b00101000000010: color_data = 12'b110011110111;
		14'b00101000000011: color_data = 12'b110011110111;
		14'b00101000000100: color_data = 12'b110011110111;
		14'b00101000000101: color_data = 12'b110011110111;
		14'b00101000000110: color_data = 12'b110011110111;
		14'b00101000000111: color_data = 12'b110011110111;
		14'b00101000001000: color_data = 12'b110011110111;
		14'b00101000001001: color_data = 12'b110011110111;
		14'b00101000001010: color_data = 12'b110011110111;
		14'b00101000001011: color_data = 12'b110011110111;
		14'b00101000001100: color_data = 12'b110011110111;
		14'b00101000001101: color_data = 12'b110011110111;
		14'b00101000001110: color_data = 12'b110011110111;
		14'b00101000001111: color_data = 12'b110011110111;
		14'b00101000010000: color_data = 12'b110011110111;
		14'b00101000010001: color_data = 12'b110011110111;
		14'b00101000010010: color_data = 12'b110011110111;
		14'b00101000010011: color_data = 12'b110011110111;
		14'b00101000011001: color_data = 12'b110011110111;
		14'b00101000011010: color_data = 12'b110011110111;
		14'b00101000011011: color_data = 12'b110011110111;
		14'b00101000011100: color_data = 12'b110011110111;
		14'b00101000011101: color_data = 12'b110011110111;
		14'b00101000100011: color_data = 12'b110011110111;
		14'b00101000100100: color_data = 12'b110011110111;
		14'b00101000100101: color_data = 12'b110011110111;
		14'b00101000100110: color_data = 12'b110011110111;
		14'b00101000100111: color_data = 12'b110011110111;
		14'b00101000101000: color_data = 12'b110011110111;
		14'b00101000101001: color_data = 12'b110011110111;
		14'b00101000101010: color_data = 12'b110011110111;
		14'b00101000101011: color_data = 12'b110011110111;
		14'b00101000101100: color_data = 12'b110011110111;
		14'b00101000101101: color_data = 12'b110011110111;
		14'b00101000101110: color_data = 12'b110011110111;
		14'b00101000101111: color_data = 12'b110011110111;
		14'b00101000110000: color_data = 12'b110011110111;
		14'b00101000110110: color_data = 12'b110011110111;
		14'b00101000110111: color_data = 12'b110011110111;
		14'b00101000111000: color_data = 12'b110011110111;
		14'b00101000111001: color_data = 12'b110011110111;
		14'b00101000111010: color_data = 12'b110011110111;
		14'b00101000111011: color_data = 12'b110011110111;
		14'b00101000111100: color_data = 12'b110011110111;
		14'b00101000111101: color_data = 12'b110011110111;
		14'b00101000111110: color_data = 12'b110011110111;
		14'b00101000111111: color_data = 12'b110011110111;
		14'b00101001000000: color_data = 12'b110011110111;
		14'b00101001000001: color_data = 12'b110011110111;
		14'b00101001000010: color_data = 12'b110011110111;
		14'b00101001000011: color_data = 12'b110011110111;
		14'b00101001000100: color_data = 12'b110011110111;
		14'b00101001001010: color_data = 12'b110011110111;
		14'b00101001001011: color_data = 12'b110011110111;
		14'b00101001001100: color_data = 12'b110011110111;
		14'b00101001001101: color_data = 12'b110011110111;
		14'b00101001001110: color_data = 12'b110011110111;
		14'b00101001010100: color_data = 12'b110011110111;
		14'b00101001010101: color_data = 12'b110011110111;
		14'b00101001010110: color_data = 12'b110011110111;
		14'b00101001010111: color_data = 12'b110011110111;
		14'b00101001011000: color_data = 12'b110011110111;
		14'b00101001011001: color_data = 12'b110011110111;
		14'b00101001011010: color_data = 12'b110011110111;
		14'b00101001011011: color_data = 12'b110011110111;
		14'b00101001011100: color_data = 12'b110011110111;
		14'b00101001011101: color_data = 12'b110011110111;
		14'b00101001011110: color_data = 12'b110011110111;
		14'b00101001011111: color_data = 12'b110011110111;
		14'b00101001100000: color_data = 12'b110011110111;
		14'b00101001100001: color_data = 12'b110011110111;
		14'b00101001101100: color_data = 12'b110011110111;
		14'b00101001101101: color_data = 12'b110011110111;
		14'b00101001101110: color_data = 12'b110011110111;
		14'b00101001101111: color_data = 12'b110011110111;
		14'b00101001110000: color_data = 12'b110011110111;
		14'b00101001110001: color_data = 12'b110011110111;
		14'b00101001110010: color_data = 12'b110011110111;
		14'b00101001110011: color_data = 12'b110011110111;
		14'b00101001110100: color_data = 12'b110011110111;
		14'b00101001110101: color_data = 12'b110011110111;
		14'b00101001110110: color_data = 12'b110011110111;
		14'b00101001110111: color_data = 12'b110011110111;
		14'b00101001111000: color_data = 12'b110011110111;
		14'b00101001111001: color_data = 12'b110011110111;
		14'b00101001111010: color_data = 12'b110011110111;
		14'b00101001111011: color_data = 12'b110011110111;
		14'b00101001111100: color_data = 12'b110011110111;
		14'b00101001111101: color_data = 12'b110011110111;
		14'b00101001111110: color_data = 12'b110011110111;
		14'b00101010000100: color_data = 12'b110011110111;
		14'b00101010000101: color_data = 12'b110011110111;
		14'b00101010000110: color_data = 12'b110011110111;
		14'b00101010000111: color_data = 12'b110011110111;
		14'b00101010001000: color_data = 12'b110011110111;
		14'b00101010010011: color_data = 12'b110011110111;
		14'b00101010010100: color_data = 12'b110011110111;
		14'b00101010010101: color_data = 12'b110011110111;
		14'b00101010010110: color_data = 12'b110011110111;
		14'b00101010010111: color_data = 12'b110011110111;
		14'b00101010011000: color_data = 12'b110011110111;
		14'b00101010011001: color_data = 12'b110011110111;
		14'b00101010011010: color_data = 12'b110011110111;
		14'b00101010011011: color_data = 12'b110011110111;
		14'b00101010011100: color_data = 12'b110011110111;
		14'b00101010100010: color_data = 12'b110011110111;
		14'b00101010100011: color_data = 12'b110011110111;
		14'b00101010100100: color_data = 12'b110011110111;
		14'b00101010100101: color_data = 12'b110011110111;
		14'b00101010100110: color_data = 12'b110011110111;
		14'b00101010101011: color_data = 12'b110011110111;
		14'b00101010101100: color_data = 12'b110011110111;
		14'b00101010101101: color_data = 12'b110011110111;
		14'b00101010101110: color_data = 12'b110011110111;
		14'b00101010101111: color_data = 12'b110011110111;
		14'b00101010110101: color_data = 12'b110011110111;
		14'b00101010110110: color_data = 12'b110011110111;
		14'b00101010110111: color_data = 12'b110011110111;
		14'b00101010111000: color_data = 12'b110011110111;
		14'b00101010111001: color_data = 12'b110011110111;
		14'b00101010111010: color_data = 12'b110011110111;
		14'b00101010111011: color_data = 12'b110011110111;
		14'b00101010111100: color_data = 12'b110011110111;
		14'b00101010111101: color_data = 12'b110011110111;
		14'b00101010111110: color_data = 12'b110011110111;
		14'b00101010111111: color_data = 12'b110011110111;
		14'b00101011000000: color_data = 12'b110011110111;
		14'b00101011000001: color_data = 12'b110011110111;
		14'b00101011000010: color_data = 12'b110011110111;
		14'b00101011000011: color_data = 12'b110011110111;
		14'b00101011001001: color_data = 12'b110011110111;
		14'b00101011001010: color_data = 12'b110011110111;
		14'b00101011001011: color_data = 12'b110011110111;
		14'b00101011001100: color_data = 12'b110011110111;
		14'b00101011001101: color_data = 12'b110011110111;
		14'b00101011001110: color_data = 12'b110011110111;
		14'b00101011001111: color_data = 12'b110011110111;
		14'b00101011010000: color_data = 12'b110011110111;
		14'b00101011010001: color_data = 12'b110011110111;
		14'b00101100000000: color_data = 12'b110011110111;
		14'b00101100000001: color_data = 12'b110011110111;
		14'b00101100000010: color_data = 12'b110011110111;
		14'b00101100000011: color_data = 12'b110011110111;
		14'b00101100000100: color_data = 12'b110011110111;
		14'b00101100000101: color_data = 12'b110011110111;
		14'b00101100000110: color_data = 12'b110011110111;
		14'b00101100000111: color_data = 12'b110011110111;
		14'b00101100001000: color_data = 12'b110011110111;
		14'b00101100001001: color_data = 12'b110011110111;
		14'b00101100001010: color_data = 12'b110011110111;
		14'b00101100001011: color_data = 12'b110011110111;
		14'b00101100001100: color_data = 12'b110011110111;
		14'b00101100001101: color_data = 12'b110011110111;
		14'b00101100001110: color_data = 12'b110011110111;
		14'b00101100001111: color_data = 12'b110011110111;
		14'b00101100010000: color_data = 12'b110011110111;
		14'b00101100010001: color_data = 12'b110011110111;
		14'b00101100010010: color_data = 12'b110011110111;
		14'b00101100010011: color_data = 12'b110011110111;
		14'b00101100011001: color_data = 12'b110011110111;
		14'b00101100011010: color_data = 12'b110011110111;
		14'b00101100011011: color_data = 12'b110011110111;
		14'b00101100011100: color_data = 12'b110011110111;
		14'b00101100011101: color_data = 12'b110011110111;
		14'b00101100100011: color_data = 12'b110011110111;
		14'b00101100100100: color_data = 12'b110011110111;
		14'b00101100100101: color_data = 12'b110011110111;
		14'b00101100100110: color_data = 12'b110011110111;
		14'b00101100100111: color_data = 12'b110011110111;
		14'b00101100101000: color_data = 12'b110011110111;
		14'b00101100101001: color_data = 12'b110011110111;
		14'b00101100101010: color_data = 12'b110011110111;
		14'b00101100101011: color_data = 12'b110011110111;
		14'b00101100101100: color_data = 12'b110011110111;
		14'b00101100101101: color_data = 12'b110011110111;
		14'b00101100101110: color_data = 12'b110011110111;
		14'b00101100101111: color_data = 12'b110011110111;
		14'b00101100110000: color_data = 12'b110011110111;
		14'b00101100110110: color_data = 12'b110011110111;
		14'b00101100110111: color_data = 12'b110011110111;
		14'b00101100111000: color_data = 12'b110011110111;
		14'b00101100111001: color_data = 12'b110011110111;
		14'b00101100111010: color_data = 12'b110011110111;
		14'b00101100111011: color_data = 12'b110011110111;
		14'b00101100111100: color_data = 12'b110011110111;
		14'b00101100111101: color_data = 12'b110011110111;
		14'b00101100111110: color_data = 12'b110011110111;
		14'b00101100111111: color_data = 12'b110011110111;
		14'b00101101000000: color_data = 12'b110011110111;
		14'b00101101000001: color_data = 12'b110011110111;
		14'b00101101000010: color_data = 12'b110011110111;
		14'b00101101000011: color_data = 12'b110011110111;
		14'b00101101000100: color_data = 12'b110011110111;
		14'b00101101001010: color_data = 12'b110011110111;
		14'b00101101001011: color_data = 12'b110011110111;
		14'b00101101001100: color_data = 12'b110011110111;
		14'b00101101001101: color_data = 12'b110011110111;
		14'b00101101001110: color_data = 12'b110011110111;
		14'b00101101010100: color_data = 12'b110011110111;
		14'b00101101010101: color_data = 12'b110011110111;
		14'b00101101010110: color_data = 12'b110011110111;
		14'b00101101010111: color_data = 12'b110011110111;
		14'b00101101011000: color_data = 12'b110011110111;
		14'b00101101011001: color_data = 12'b110011110111;
		14'b00101101011010: color_data = 12'b110011110111;
		14'b00101101011011: color_data = 12'b110011110111;
		14'b00101101011100: color_data = 12'b110011110111;
		14'b00101101011101: color_data = 12'b110011110111;
		14'b00101101011110: color_data = 12'b110011110111;
		14'b00101101011111: color_data = 12'b110011110111;
		14'b00101101100000: color_data = 12'b110011110111;
		14'b00101101100001: color_data = 12'b110011110111;
		14'b00101101101100: color_data = 12'b110011110111;
		14'b00101101101101: color_data = 12'b110011110111;
		14'b00101101101110: color_data = 12'b110011110111;
		14'b00101101101111: color_data = 12'b110011110111;
		14'b00101101110000: color_data = 12'b110011110111;
		14'b00101101110001: color_data = 12'b110011110111;
		14'b00101101110010: color_data = 12'b110011110111;
		14'b00101101110011: color_data = 12'b110011110111;
		14'b00101101110100: color_data = 12'b110011110111;
		14'b00101101110101: color_data = 12'b110011110111;
		14'b00101101110110: color_data = 12'b110011110111;
		14'b00101101110111: color_data = 12'b110011110111;
		14'b00101101111000: color_data = 12'b110011110111;
		14'b00101101111001: color_data = 12'b110011110111;
		14'b00101101111010: color_data = 12'b110011110111;
		14'b00101101111011: color_data = 12'b110011110111;
		14'b00101101111100: color_data = 12'b110011110111;
		14'b00101101111101: color_data = 12'b110011110111;
		14'b00101101111110: color_data = 12'b110011110111;
		14'b00101110000100: color_data = 12'b110011110111;
		14'b00101110000101: color_data = 12'b110011110111;
		14'b00101110000110: color_data = 12'b110011110111;
		14'b00101110000111: color_data = 12'b110011110111;
		14'b00101110001000: color_data = 12'b110011110111;
		14'b00101110010011: color_data = 12'b110011110111;
		14'b00101110010100: color_data = 12'b110011110111;
		14'b00101110010101: color_data = 12'b110011110111;
		14'b00101110010110: color_data = 12'b110011110111;
		14'b00101110010111: color_data = 12'b110011110111;
		14'b00101110011000: color_data = 12'b110011110111;
		14'b00101110011001: color_data = 12'b110011110111;
		14'b00101110011010: color_data = 12'b110011110111;
		14'b00101110011011: color_data = 12'b110011110111;
		14'b00101110011100: color_data = 12'b110011110111;
		14'b00101110100010: color_data = 12'b110011110111;
		14'b00101110100011: color_data = 12'b110011110111;
		14'b00101110100100: color_data = 12'b110011110111;
		14'b00101110100101: color_data = 12'b110011110111;
		14'b00101110100110: color_data = 12'b110011110111;
		14'b00101110101011: color_data = 12'b110011110111;
		14'b00101110101100: color_data = 12'b110011110111;
		14'b00101110101101: color_data = 12'b110011110111;
		14'b00101110101110: color_data = 12'b110011110111;
		14'b00101110101111: color_data = 12'b110011110111;
		14'b00101110110101: color_data = 12'b110011110111;
		14'b00101110110110: color_data = 12'b110011110111;
		14'b00101110110111: color_data = 12'b110011110111;
		14'b00101110111000: color_data = 12'b110011110111;
		14'b00101110111001: color_data = 12'b110011110111;
		14'b00101110111010: color_data = 12'b110011110111;
		14'b00101110111011: color_data = 12'b110011110111;
		14'b00101110111100: color_data = 12'b110011110111;
		14'b00101110111101: color_data = 12'b110011110111;
		14'b00101110111110: color_data = 12'b110011110111;
		14'b00101110111111: color_data = 12'b110011110111;
		14'b00101111000000: color_data = 12'b110011110111;
		14'b00101111000001: color_data = 12'b110011110111;
		14'b00101111000010: color_data = 12'b110011110111;
		14'b00101111000011: color_data = 12'b110011110111;
		14'b00101111001001: color_data = 12'b110011110111;
		14'b00101111001010: color_data = 12'b110011110111;
		14'b00101111001011: color_data = 12'b110011110111;
		14'b00101111001100: color_data = 12'b110011110111;
		14'b00101111001101: color_data = 12'b110011110111;
		14'b00101111001110: color_data = 12'b110011110111;
		14'b00101111001111: color_data = 12'b110011110111;
		14'b00101111010000: color_data = 12'b110011110111;
		14'b00101111010001: color_data = 12'b110011110111;
		14'b00110000000000: color_data = 12'b110011110111;
		14'b00110000000001: color_data = 12'b110011110111;
		14'b00110000000010: color_data = 12'b110011110111;
		14'b00110000000011: color_data = 12'b110011110111;
		14'b00110000000100: color_data = 12'b110011110111;
		14'b00110000000101: color_data = 12'b110011110111;
		14'b00110000000110: color_data = 12'b110011110111;
		14'b00110000000111: color_data = 12'b110011110111;
		14'b00110000001000: color_data = 12'b110011110111;
		14'b00110000001001: color_data = 12'b110011110111;
		14'b00110000001010: color_data = 12'b110011110111;
		14'b00110000001011: color_data = 12'b110011110111;
		14'b00110000001100: color_data = 12'b110011110111;
		14'b00110000001101: color_data = 12'b110011110111;
		14'b00110000001110: color_data = 12'b110011110111;
		14'b00110000001111: color_data = 12'b110011110111;
		14'b00110000010000: color_data = 12'b110011110111;
		14'b00110000010001: color_data = 12'b110011110111;
		14'b00110000010010: color_data = 12'b110011110111;
		14'b00110000010011: color_data = 12'b110011110111;
		14'b00110000011001: color_data = 12'b110011110111;
		14'b00110000011010: color_data = 12'b110011110111;
		14'b00110000011011: color_data = 12'b110011110111;
		14'b00110000011100: color_data = 12'b110011110111;
		14'b00110000011101: color_data = 12'b110011110111;
		14'b00110000100011: color_data = 12'b110011110111;
		14'b00110000100100: color_data = 12'b110011110111;
		14'b00110000100101: color_data = 12'b110011110111;
		14'b00110000100110: color_data = 12'b110011110111;
		14'b00110000100111: color_data = 12'b110011110111;
		14'b00110000101000: color_data = 12'b110011110111;
		14'b00110000101001: color_data = 12'b110011110111;
		14'b00110000101010: color_data = 12'b110011110111;
		14'b00110000101011: color_data = 12'b110011110111;
		14'b00110000101100: color_data = 12'b110011110111;
		14'b00110000101101: color_data = 12'b110011110111;
		14'b00110000101110: color_data = 12'b110011110111;
		14'b00110000101111: color_data = 12'b110011110111;
		14'b00110000110000: color_data = 12'b110011110111;
		14'b00110000110110: color_data = 12'b110011110111;
		14'b00110000110111: color_data = 12'b110011110111;
		14'b00110000111000: color_data = 12'b110011110111;
		14'b00110000111001: color_data = 12'b110011110111;
		14'b00110000111010: color_data = 12'b110011110111;
		14'b00110000111011: color_data = 12'b110011110111;
		14'b00110000111100: color_data = 12'b110011110111;
		14'b00110000111101: color_data = 12'b110011110111;
		14'b00110000111110: color_data = 12'b110011110111;
		14'b00110000111111: color_data = 12'b110011110111;
		14'b00110001000000: color_data = 12'b110011110111;
		14'b00110001000001: color_data = 12'b110011110111;
		14'b00110001000010: color_data = 12'b110011110111;
		14'b00110001000011: color_data = 12'b110011110111;
		14'b00110001000100: color_data = 12'b110011110111;
		14'b00110001001010: color_data = 12'b110011110111;
		14'b00110001001011: color_data = 12'b110011110111;
		14'b00110001001100: color_data = 12'b110011110111;
		14'b00110001001101: color_data = 12'b110011110111;
		14'b00110001001110: color_data = 12'b110011110111;
		14'b00110001010100: color_data = 12'b110011110111;
		14'b00110001010101: color_data = 12'b110011110111;
		14'b00110001010110: color_data = 12'b110011110111;
		14'b00110001010111: color_data = 12'b110011110111;
		14'b00110001011000: color_data = 12'b110011110111;
		14'b00110001011001: color_data = 12'b110011110111;
		14'b00110001011010: color_data = 12'b110011110111;
		14'b00110001011011: color_data = 12'b110011110111;
		14'b00110001011100: color_data = 12'b110011110111;
		14'b00110001011101: color_data = 12'b110011110111;
		14'b00110001011110: color_data = 12'b110011110111;
		14'b00110001011111: color_data = 12'b110011110111;
		14'b00110001100000: color_data = 12'b110011110111;
		14'b00110001100001: color_data = 12'b110011110111;
		14'b00110001101100: color_data = 12'b110011110111;
		14'b00110001101101: color_data = 12'b110011110111;
		14'b00110001101110: color_data = 12'b110011110111;
		14'b00110001101111: color_data = 12'b110011110111;
		14'b00110001110000: color_data = 12'b110011110111;
		14'b00110001110001: color_data = 12'b110011110111;
		14'b00110001110010: color_data = 12'b110011110111;
		14'b00110001110011: color_data = 12'b110011110111;
		14'b00110001110100: color_data = 12'b110011110111;
		14'b00110001110101: color_data = 12'b110011110111;
		14'b00110001110110: color_data = 12'b110011110111;
		14'b00110001110111: color_data = 12'b110011110111;
		14'b00110001111000: color_data = 12'b110011110111;
		14'b00110001111001: color_data = 12'b110011110111;
		14'b00110001111010: color_data = 12'b110011110111;
		14'b00110001111011: color_data = 12'b110011110111;
		14'b00110001111100: color_data = 12'b110011110111;
		14'b00110001111101: color_data = 12'b110011110111;
		14'b00110001111110: color_data = 12'b110011110111;
		14'b00110010000100: color_data = 12'b110011110111;
		14'b00110010000101: color_data = 12'b110011110111;
		14'b00110010000110: color_data = 12'b110011110111;
		14'b00110010000111: color_data = 12'b110011110111;
		14'b00110010001000: color_data = 12'b110011110111;
		14'b00110010010011: color_data = 12'b110011110111;
		14'b00110010010100: color_data = 12'b110011110111;
		14'b00110010010101: color_data = 12'b110011110111;
		14'b00110010010110: color_data = 12'b110011110111;
		14'b00110010010111: color_data = 12'b110011110111;
		14'b00110010011000: color_data = 12'b110011110111;
		14'b00110010011001: color_data = 12'b110011110111;
		14'b00110010011010: color_data = 12'b110011110111;
		14'b00110010011011: color_data = 12'b110011110111;
		14'b00110010011100: color_data = 12'b110011110111;
		14'b00110010100010: color_data = 12'b110011110111;
		14'b00110010100011: color_data = 12'b110011110111;
		14'b00110010100100: color_data = 12'b110011110111;
		14'b00110010100101: color_data = 12'b110011110111;
		14'b00110010100110: color_data = 12'b110011110111;
		14'b00110010101011: color_data = 12'b110011110111;
		14'b00110010101100: color_data = 12'b110011110111;
		14'b00110010101101: color_data = 12'b110011110111;
		14'b00110010101110: color_data = 12'b110011110111;
		14'b00110010101111: color_data = 12'b110011110111;
		14'b00110010110101: color_data = 12'b110011110111;
		14'b00110010110110: color_data = 12'b110011110111;
		14'b00110010110111: color_data = 12'b110011110111;
		14'b00110010111000: color_data = 12'b110011110111;
		14'b00110010111001: color_data = 12'b110011110111;
		14'b00110010111010: color_data = 12'b110011110111;
		14'b00110010111011: color_data = 12'b110011110111;
		14'b00110010111100: color_data = 12'b110011110111;
		14'b00110010111101: color_data = 12'b110011110111;
		14'b00110010111110: color_data = 12'b110011110111;
		14'b00110010111111: color_data = 12'b110011110111;
		14'b00110011000000: color_data = 12'b110011110111;
		14'b00110011000001: color_data = 12'b110011110111;
		14'b00110011000010: color_data = 12'b110011110111;
		14'b00110011000011: color_data = 12'b110011110111;
		14'b00110011001001: color_data = 12'b110011110111;
		14'b00110011001010: color_data = 12'b110011110111;
		14'b00110011001011: color_data = 12'b110011110111;
		14'b00110011001100: color_data = 12'b110011110111;
		14'b00110011001101: color_data = 12'b110011110111;
		14'b00110011001110: color_data = 12'b110011110111;
		14'b00110011001111: color_data = 12'b110011110111;
		14'b00110011010000: color_data = 12'b110011110111;
		14'b00110011010001: color_data = 12'b110011110111;
		14'b00110100000000: color_data = 12'b110011110111;
		14'b00110100000001: color_data = 12'b110011110111;
		14'b00110100000010: color_data = 12'b110011110111;
		14'b00110100000011: color_data = 12'b110011110111;
		14'b00110100000100: color_data = 12'b110011110111;
		14'b00110100000101: color_data = 12'b110011110111;
		14'b00110100000110: color_data = 12'b110011110111;
		14'b00110100000111: color_data = 12'b110011110111;
		14'b00110100001000: color_data = 12'b110011110111;
		14'b00110100001001: color_data = 12'b110011110111;
		14'b00110100001010: color_data = 12'b110011110111;
		14'b00110100001011: color_data = 12'b110011110111;
		14'b00110100001100: color_data = 12'b110011110111;
		14'b00110100001101: color_data = 12'b110011110111;
		14'b00110100001110: color_data = 12'b110011110111;
		14'b00110100001111: color_data = 12'b110011110111;
		14'b00110100010000: color_data = 12'b110011110111;
		14'b00110100010001: color_data = 12'b110011110111;
		14'b00110100010010: color_data = 12'b110011110111;
		14'b00110100010011: color_data = 12'b110011110111;
		14'b00110100011001: color_data = 12'b110011110111;
		14'b00110100011010: color_data = 12'b110011110111;
		14'b00110100011011: color_data = 12'b110011110111;
		14'b00110100011100: color_data = 12'b110011110111;
		14'b00110100011101: color_data = 12'b110011110111;
		14'b00110100100011: color_data = 12'b110011110111;
		14'b00110100100100: color_data = 12'b110011110111;
		14'b00110100100101: color_data = 12'b110011110111;
		14'b00110100100110: color_data = 12'b110011110111;
		14'b00110100100111: color_data = 12'b110011110111;
		14'b00110100101000: color_data = 12'b110011110111;
		14'b00110100101001: color_data = 12'b110011110111;
		14'b00110100101010: color_data = 12'b110011110111;
		14'b00110100101011: color_data = 12'b110011110111;
		14'b00110100101100: color_data = 12'b110011110111;
		14'b00110100101101: color_data = 12'b110011110111;
		14'b00110100101110: color_data = 12'b110011110111;
		14'b00110100101111: color_data = 12'b110011110111;
		14'b00110100110000: color_data = 12'b110011110111;
		14'b00110100110110: color_data = 12'b110011110111;
		14'b00110100110111: color_data = 12'b110011110111;
		14'b00110100111000: color_data = 12'b110011110111;
		14'b00110100111001: color_data = 12'b110011110111;
		14'b00110100111010: color_data = 12'b110011110111;
		14'b00110100111011: color_data = 12'b110011110111;
		14'b00110100111100: color_data = 12'b110011110111;
		14'b00110100111101: color_data = 12'b110011110111;
		14'b00110100111110: color_data = 12'b110011110111;
		14'b00110100111111: color_data = 12'b110011110111;
		14'b00110101000000: color_data = 12'b110011110111;
		14'b00110101000001: color_data = 12'b110011110111;
		14'b00110101000010: color_data = 12'b110011110111;
		14'b00110101000011: color_data = 12'b110011110111;
		14'b00110101000100: color_data = 12'b110011110111;
		14'b00110101001010: color_data = 12'b110011110111;
		14'b00110101001011: color_data = 12'b110011110111;
		14'b00110101001100: color_data = 12'b110011110111;
		14'b00110101001101: color_data = 12'b110011110111;
		14'b00110101001110: color_data = 12'b110011110111;
		14'b00110101010100: color_data = 12'b110011110111;
		14'b00110101010101: color_data = 12'b110011110111;
		14'b00110101010110: color_data = 12'b110011110111;
		14'b00110101010111: color_data = 12'b110011110111;
		14'b00110101011000: color_data = 12'b110011110111;
		14'b00110101011001: color_data = 12'b110011110111;
		14'b00110101011010: color_data = 12'b110011110111;
		14'b00110101011011: color_data = 12'b110011110111;
		14'b00110101011100: color_data = 12'b110011110111;
		14'b00110101011101: color_data = 12'b110011110111;
		14'b00110101011110: color_data = 12'b110011110111;
		14'b00110101011111: color_data = 12'b110011110111;
		14'b00110101100000: color_data = 12'b110011110111;
		14'b00110101100001: color_data = 12'b110011110111;
		14'b00110101101100: color_data = 12'b110011110111;
		14'b00110101101101: color_data = 12'b110011110111;
		14'b00110101101110: color_data = 12'b110011110111;
		14'b00110101101111: color_data = 12'b110011110111;
		14'b00110101110000: color_data = 12'b110011110111;
		14'b00110101110001: color_data = 12'b110011110111;
		14'b00110101110010: color_data = 12'b110011110111;
		14'b00110101110011: color_data = 12'b110011110111;
		14'b00110101110100: color_data = 12'b110011110111;
		14'b00110101110101: color_data = 12'b110011110111;
		14'b00110101110110: color_data = 12'b110011110111;
		14'b00110101110111: color_data = 12'b110011110111;
		14'b00110101111000: color_data = 12'b110011110111;
		14'b00110101111001: color_data = 12'b110011110111;
		14'b00110101111010: color_data = 12'b110011110111;
		14'b00110101111011: color_data = 12'b110011110111;
		14'b00110101111100: color_data = 12'b110011110111;
		14'b00110101111101: color_data = 12'b110011110111;
		14'b00110101111110: color_data = 12'b110011110111;
		14'b00110110000100: color_data = 12'b110011110111;
		14'b00110110000101: color_data = 12'b110011110111;
		14'b00110110000110: color_data = 12'b110011110111;
		14'b00110110000111: color_data = 12'b110011110111;
		14'b00110110001000: color_data = 12'b110011110111;
		14'b00110110010011: color_data = 12'b110011110111;
		14'b00110110010100: color_data = 12'b110011110111;
		14'b00110110010101: color_data = 12'b110011110111;
		14'b00110110010110: color_data = 12'b110011110111;
		14'b00110110010111: color_data = 12'b110011110111;
		14'b00110110011000: color_data = 12'b110011110111;
		14'b00110110011001: color_data = 12'b110011110111;
		14'b00110110011010: color_data = 12'b110011110111;
		14'b00110110011011: color_data = 12'b110011110111;
		14'b00110110011100: color_data = 12'b110011110111;
		14'b00110110100010: color_data = 12'b110011110111;
		14'b00110110100011: color_data = 12'b110011110111;
		14'b00110110100100: color_data = 12'b110011110111;
		14'b00110110100101: color_data = 12'b110011110111;
		14'b00110110100110: color_data = 12'b110011110111;
		14'b00110110101011: color_data = 12'b110011110111;
		14'b00110110101100: color_data = 12'b110011110111;
		14'b00110110101101: color_data = 12'b110011110111;
		14'b00110110101110: color_data = 12'b110011110111;
		14'b00110110101111: color_data = 12'b110011110111;
		14'b00110110110101: color_data = 12'b110011110111;
		14'b00110110110110: color_data = 12'b110011110111;
		14'b00110110110111: color_data = 12'b110011110111;
		14'b00110110111000: color_data = 12'b110011110111;
		14'b00110110111001: color_data = 12'b110011110111;
		14'b00110110111010: color_data = 12'b110011110111;
		14'b00110110111011: color_data = 12'b110011110111;
		14'b00110110111100: color_data = 12'b110011110111;
		14'b00110110111101: color_data = 12'b110011110111;
		14'b00110110111110: color_data = 12'b110011110111;
		14'b00110110111111: color_data = 12'b110011110111;
		14'b00110111000000: color_data = 12'b110011110111;
		14'b00110111000001: color_data = 12'b110011110111;
		14'b00110111000010: color_data = 12'b110011110111;
		14'b00110111000011: color_data = 12'b110011110111;
		14'b00110111001001: color_data = 12'b110011110111;
		14'b00110111001010: color_data = 12'b110011110111;
		14'b00110111001011: color_data = 12'b110011110111;
		14'b00110111001100: color_data = 12'b110011110111;
		14'b00110111001101: color_data = 12'b110011110111;
		14'b00110111001110: color_data = 12'b110011110111;
		14'b00110111001111: color_data = 12'b110011110111;
		14'b00110111010000: color_data = 12'b110011110111;
		14'b00110111010001: color_data = 12'b110011110111;
		14'b00111000001111: color_data = 12'b110011110111;
		14'b00111000010000: color_data = 12'b110011110111;
		14'b00111000010001: color_data = 12'b110011110111;
		14'b00111000010010: color_data = 12'b110011110111;
		14'b00111000010011: color_data = 12'b110011110111;
		14'b00111000011001: color_data = 12'b110011110111;
		14'b00111000011010: color_data = 12'b110011110111;
		14'b00111000011011: color_data = 12'b110011110111;
		14'b00111000011100: color_data = 12'b110011110111;
		14'b00111000011101: color_data = 12'b110011110111;
		14'b00111000100011: color_data = 12'b110011110111;
		14'b00111000100100: color_data = 12'b110011110111;
		14'b00111000100101: color_data = 12'b110011110111;
		14'b00111000100110: color_data = 12'b110011110111;
		14'b00111000100111: color_data = 12'b110011110111;
		14'b00111000101100: color_data = 12'b110011110111;
		14'b00111000101101: color_data = 12'b110011110111;
		14'b00111000101110: color_data = 12'b110011110111;
		14'b00111000101111: color_data = 12'b110011110111;
		14'b00111000110000: color_data = 12'b110011110111;
		14'b00111000110110: color_data = 12'b110011110111;
		14'b00111000110111: color_data = 12'b110011110111;
		14'b00111000111000: color_data = 12'b110011110111;
		14'b00111000111001: color_data = 12'b110011110111;
		14'b00111000111010: color_data = 12'b110011110111;
		14'b00111001000000: color_data = 12'b110011110111;
		14'b00111001000001: color_data = 12'b110011110111;
		14'b00111001000010: color_data = 12'b110011110111;
		14'b00111001000011: color_data = 12'b110011110111;
		14'b00111001000100: color_data = 12'b110011110111;
		14'b00111001001010: color_data = 12'b110011110111;
		14'b00111001001011: color_data = 12'b110011110111;
		14'b00111001001100: color_data = 12'b110011110111;
		14'b00111001001101: color_data = 12'b110011110111;
		14'b00111001001110: color_data = 12'b110011110111;
		14'b00111001010100: color_data = 12'b110011110111;
		14'b00111001010101: color_data = 12'b110011110111;
		14'b00111001010110: color_data = 12'b110011110111;
		14'b00111001010111: color_data = 12'b110011110111;
		14'b00111001011101: color_data = 12'b110011110111;
		14'b00111001011110: color_data = 12'b110011110111;
		14'b00111001011111: color_data = 12'b110011110111;
		14'b00111001100000: color_data = 12'b110011110111;
		14'b00111001100001: color_data = 12'b110011110111;
		14'b00111001101100: color_data = 12'b110011110111;
		14'b00111001101101: color_data = 12'b110011110111;
		14'b00111001101110: color_data = 12'b110011110111;
		14'b00111001101111: color_data = 12'b110011110111;
		14'b00111001110000: color_data = 12'b110011110111;
		14'b00111010000100: color_data = 12'b110011110111;
		14'b00111010000101: color_data = 12'b110011110111;
		14'b00111010000110: color_data = 12'b110011110111;
		14'b00111010000111: color_data = 12'b110011110111;
		14'b00111010001000: color_data = 12'b110011110111;
		14'b00111010001110: color_data = 12'b110011110111;
		14'b00111010001111: color_data = 12'b110011110111;
		14'b00111010010000: color_data = 12'b110011110111;
		14'b00111010010001: color_data = 12'b110011110111;
		14'b00111010010010: color_data = 12'b110011110111;
		14'b00111010011000: color_data = 12'b110011110111;
		14'b00111010011001: color_data = 12'b110011110111;
		14'b00111010011010: color_data = 12'b110011110111;
		14'b00111010011011: color_data = 12'b110011110111;
		14'b00111010011100: color_data = 12'b110011110111;
		14'b00111010100010: color_data = 12'b110011110111;
		14'b00111010100011: color_data = 12'b110011110111;
		14'b00111010100100: color_data = 12'b110011110111;
		14'b00111010100101: color_data = 12'b110011110111;
		14'b00111010100110: color_data = 12'b110011110111;
		14'b00111010101011: color_data = 12'b110011110111;
		14'b00111010101100: color_data = 12'b110011110111;
		14'b00111010101101: color_data = 12'b110011110111;
		14'b00111010101110: color_data = 12'b110011110111;
		14'b00111010101111: color_data = 12'b110011110111;
		14'b00111010110101: color_data = 12'b110011110111;
		14'b00111010110110: color_data = 12'b110011110111;
		14'b00111010110111: color_data = 12'b110011110111;
		14'b00111010111000: color_data = 12'b110011110111;
		14'b00111010111001: color_data = 12'b110011110111;
		14'b00111010111111: color_data = 12'b110011110111;
		14'b00111011000000: color_data = 12'b110011110111;
		14'b00111011000001: color_data = 12'b110011110111;
		14'b00111011000010: color_data = 12'b110011110111;
		14'b00111011000011: color_data = 12'b110011110111;
		14'b00111011001001: color_data = 12'b110011110111;
		14'b00111011001010: color_data = 12'b110011110111;
		14'b00111011001011: color_data = 12'b110011110111;
		14'b00111011001100: color_data = 12'b110011110111;
		14'b00111011001101: color_data = 12'b110011110111;
		14'b00111100001111: color_data = 12'b110011110111;
		14'b00111100010000: color_data = 12'b110011110111;
		14'b00111100010001: color_data = 12'b110011110111;
		14'b00111100010010: color_data = 12'b110011110111;
		14'b00111100010011: color_data = 12'b110011110111;
		14'b00111100011001: color_data = 12'b110011110111;
		14'b00111100011010: color_data = 12'b110011110111;
		14'b00111100011011: color_data = 12'b110011110111;
		14'b00111100011100: color_data = 12'b110011110111;
		14'b00111100011101: color_data = 12'b110011110111;
		14'b00111100100011: color_data = 12'b110011110111;
		14'b00111100100100: color_data = 12'b110011110111;
		14'b00111100100101: color_data = 12'b110011110111;
		14'b00111100100110: color_data = 12'b110011110111;
		14'b00111100100111: color_data = 12'b110011110111;
		14'b00111100101100: color_data = 12'b110011110111;
		14'b00111100101101: color_data = 12'b110011110111;
		14'b00111100101110: color_data = 12'b110011110111;
		14'b00111100101111: color_data = 12'b110011110111;
		14'b00111100110000: color_data = 12'b110011110111;
		14'b00111100110110: color_data = 12'b110011110111;
		14'b00111100110111: color_data = 12'b110011110111;
		14'b00111100111000: color_data = 12'b110011110111;
		14'b00111100111001: color_data = 12'b110011110111;
		14'b00111100111010: color_data = 12'b110011110111;
		14'b00111101000000: color_data = 12'b110011110111;
		14'b00111101000001: color_data = 12'b110011110111;
		14'b00111101000010: color_data = 12'b110011110111;
		14'b00111101000011: color_data = 12'b110011110111;
		14'b00111101000100: color_data = 12'b110011110111;
		14'b00111101001010: color_data = 12'b110011110111;
		14'b00111101001011: color_data = 12'b110011110111;
		14'b00111101001100: color_data = 12'b110011110111;
		14'b00111101001101: color_data = 12'b110011110111;
		14'b00111101001110: color_data = 12'b110011110111;
		14'b00111101010100: color_data = 12'b110011110111;
		14'b00111101010101: color_data = 12'b110011110111;
		14'b00111101010110: color_data = 12'b110011110111;
		14'b00111101010111: color_data = 12'b110011110111;
		14'b00111101011101: color_data = 12'b110011110111;
		14'b00111101011110: color_data = 12'b110011110111;
		14'b00111101011111: color_data = 12'b110011110111;
		14'b00111101100000: color_data = 12'b110011110111;
		14'b00111101100001: color_data = 12'b110011110111;
		14'b00111101101100: color_data = 12'b110011110111;
		14'b00111101101101: color_data = 12'b110011110111;
		14'b00111101101110: color_data = 12'b110011110111;
		14'b00111101101111: color_data = 12'b110011110111;
		14'b00111101110000: color_data = 12'b110011110111;
		14'b00111110000100: color_data = 12'b110011110111;
		14'b00111110000101: color_data = 12'b110011110111;
		14'b00111110000110: color_data = 12'b110011110111;
		14'b00111110000111: color_data = 12'b110011110111;
		14'b00111110001000: color_data = 12'b110011110111;
		14'b00111110001110: color_data = 12'b110011110111;
		14'b00111110001111: color_data = 12'b110011110111;
		14'b00111110010000: color_data = 12'b110011110111;
		14'b00111110010001: color_data = 12'b110011110111;
		14'b00111110010010: color_data = 12'b110011110111;
		14'b00111110011000: color_data = 12'b110011110111;
		14'b00111110011001: color_data = 12'b110011110111;
		14'b00111110011010: color_data = 12'b110011110111;
		14'b00111110011011: color_data = 12'b110011110111;
		14'b00111110011100: color_data = 12'b110011110111;
		14'b00111110100010: color_data = 12'b110011110111;
		14'b00111110100011: color_data = 12'b110011110111;
		14'b00111110100100: color_data = 12'b110011110111;
		14'b00111110100101: color_data = 12'b110011110111;
		14'b00111110100110: color_data = 12'b110011110111;
		14'b00111110101011: color_data = 12'b110011110111;
		14'b00111110101100: color_data = 12'b110011110111;
		14'b00111110101101: color_data = 12'b110011110111;
		14'b00111110101110: color_data = 12'b110011110111;
		14'b00111110101111: color_data = 12'b110011110111;
		14'b00111110110101: color_data = 12'b110011110111;
		14'b00111110110110: color_data = 12'b110011110111;
		14'b00111110110111: color_data = 12'b110011110111;
		14'b00111110111000: color_data = 12'b110011110111;
		14'b00111110111001: color_data = 12'b110011110111;
		14'b00111110111111: color_data = 12'b110011110111;
		14'b00111111000000: color_data = 12'b110011110111;
		14'b00111111000001: color_data = 12'b110011110111;
		14'b00111111000010: color_data = 12'b110011110111;
		14'b00111111000011: color_data = 12'b110011110111;
		14'b00111111001001: color_data = 12'b110011110111;
		14'b00111111001010: color_data = 12'b110011110111;
		14'b00111111001011: color_data = 12'b110011110111;
		14'b00111111001100: color_data = 12'b110011110111;
		14'b00111111001101: color_data = 12'b110011110111;
		14'b01000000001111: color_data = 12'b110011110111;
		14'b01000000010000: color_data = 12'b110011110111;
		14'b01000000010001: color_data = 12'b110011110111;
		14'b01000000010010: color_data = 12'b110011110111;
		14'b01000000010011: color_data = 12'b110011110111;
		14'b01000000011001: color_data = 12'b110011110111;
		14'b01000000011010: color_data = 12'b110011110111;
		14'b01000000011011: color_data = 12'b110011110111;
		14'b01000000011100: color_data = 12'b110011110111;
		14'b01000000011101: color_data = 12'b110011110111;
		14'b01000000100011: color_data = 12'b110011110111;
		14'b01000000100100: color_data = 12'b110011110111;
		14'b01000000100101: color_data = 12'b110011110111;
		14'b01000000100110: color_data = 12'b110011110111;
		14'b01000000100111: color_data = 12'b110011110111;
		14'b01000000101100: color_data = 12'b110011110111;
		14'b01000000101101: color_data = 12'b110011110111;
		14'b01000000101110: color_data = 12'b110011110111;
		14'b01000000101111: color_data = 12'b110011110111;
		14'b01000000110000: color_data = 12'b110011110111;
		14'b01000000110110: color_data = 12'b110011110111;
		14'b01000000110111: color_data = 12'b110011110111;
		14'b01000000111000: color_data = 12'b110011110111;
		14'b01000000111001: color_data = 12'b110011110111;
		14'b01000000111010: color_data = 12'b110011110111;
		14'b01000001000000: color_data = 12'b110011110111;
		14'b01000001000001: color_data = 12'b110011110111;
		14'b01000001000010: color_data = 12'b110011110111;
		14'b01000001000011: color_data = 12'b110011110111;
		14'b01000001000100: color_data = 12'b110011110111;
		14'b01000001001010: color_data = 12'b110011110111;
		14'b01000001001011: color_data = 12'b110011110111;
		14'b01000001001100: color_data = 12'b110011110111;
		14'b01000001001101: color_data = 12'b110011110111;
		14'b01000001001110: color_data = 12'b110011110111;
		14'b01000001010100: color_data = 12'b110011110111;
		14'b01000001010101: color_data = 12'b110011110111;
		14'b01000001010110: color_data = 12'b110011110111;
		14'b01000001010111: color_data = 12'b110011110111;
		14'b01000001011101: color_data = 12'b110011110111;
		14'b01000001011110: color_data = 12'b110011110111;
		14'b01000001011111: color_data = 12'b110011110111;
		14'b01000001100000: color_data = 12'b110011110111;
		14'b01000001100001: color_data = 12'b110011110111;
		14'b01000001101100: color_data = 12'b110011110111;
		14'b01000001101101: color_data = 12'b110011110111;
		14'b01000001101110: color_data = 12'b110011110111;
		14'b01000001101111: color_data = 12'b110011110111;
		14'b01000001110000: color_data = 12'b110011110111;
		14'b01000010000100: color_data = 12'b110011110111;
		14'b01000010000101: color_data = 12'b110011110111;
		14'b01000010000110: color_data = 12'b110011110111;
		14'b01000010000111: color_data = 12'b110011110111;
		14'b01000010001000: color_data = 12'b110011110111;
		14'b01000010001110: color_data = 12'b110011110111;
		14'b01000010001111: color_data = 12'b110011110111;
		14'b01000010010000: color_data = 12'b110011110111;
		14'b01000010010001: color_data = 12'b110011110111;
		14'b01000010010010: color_data = 12'b110011110111;
		14'b01000010011000: color_data = 12'b110011110111;
		14'b01000010011001: color_data = 12'b110011110111;
		14'b01000010011010: color_data = 12'b110011110111;
		14'b01000010011011: color_data = 12'b110011110111;
		14'b01000010011100: color_data = 12'b110011110111;
		14'b01000010100010: color_data = 12'b110011110111;
		14'b01000010100011: color_data = 12'b110011110111;
		14'b01000010100100: color_data = 12'b110011110111;
		14'b01000010100101: color_data = 12'b110011110111;
		14'b01000010100110: color_data = 12'b110011110111;
		14'b01000010101011: color_data = 12'b110011110111;
		14'b01000010101100: color_data = 12'b110011110111;
		14'b01000010101101: color_data = 12'b110011110111;
		14'b01000010101110: color_data = 12'b110011110111;
		14'b01000010101111: color_data = 12'b110011110111;
		14'b01000010110101: color_data = 12'b110011110111;
		14'b01000010110110: color_data = 12'b110011110111;
		14'b01000010110111: color_data = 12'b110011110111;
		14'b01000010111000: color_data = 12'b110011110111;
		14'b01000010111001: color_data = 12'b110011110111;
		14'b01000010111111: color_data = 12'b110011110111;
		14'b01000011000000: color_data = 12'b110011110111;
		14'b01000011000001: color_data = 12'b110011110111;
		14'b01000011000010: color_data = 12'b110011110111;
		14'b01000011000011: color_data = 12'b110011110111;
		14'b01000011001001: color_data = 12'b110011110111;
		14'b01000011001010: color_data = 12'b110011110111;
		14'b01000011001011: color_data = 12'b110011110111;
		14'b01000011001100: color_data = 12'b110011110111;
		14'b01000011001101: color_data = 12'b110011110111;
		14'b01000100001111: color_data = 12'b110011110111;
		14'b01000100010000: color_data = 12'b110011110111;
		14'b01000100010001: color_data = 12'b110011110111;
		14'b01000100010010: color_data = 12'b110011110111;
		14'b01000100010011: color_data = 12'b110011110111;
		14'b01000100011001: color_data = 12'b110011110111;
		14'b01000100011010: color_data = 12'b110011110111;
		14'b01000100011011: color_data = 12'b110011110111;
		14'b01000100011100: color_data = 12'b110011110111;
		14'b01000100011101: color_data = 12'b110011110111;
		14'b01000100100011: color_data = 12'b110011110111;
		14'b01000100100100: color_data = 12'b110011110111;
		14'b01000100100101: color_data = 12'b110011110111;
		14'b01000100100110: color_data = 12'b110011110111;
		14'b01000100100111: color_data = 12'b110011110111;
		14'b01000100101100: color_data = 12'b110011110111;
		14'b01000100101101: color_data = 12'b110011110111;
		14'b01000100101110: color_data = 12'b110011110111;
		14'b01000100101111: color_data = 12'b110011110111;
		14'b01000100110000: color_data = 12'b110011110111;
		14'b01000100110110: color_data = 12'b110011110111;
		14'b01000100110111: color_data = 12'b110011110111;
		14'b01000100111000: color_data = 12'b110011110111;
		14'b01000100111001: color_data = 12'b110011110111;
		14'b01000100111010: color_data = 12'b110011110111;
		14'b01000101000000: color_data = 12'b110011110111;
		14'b01000101000001: color_data = 12'b110011110111;
		14'b01000101000010: color_data = 12'b110011110111;
		14'b01000101000011: color_data = 12'b110011110111;
		14'b01000101000100: color_data = 12'b110011110111;
		14'b01000101001010: color_data = 12'b110011110111;
		14'b01000101001011: color_data = 12'b110011110111;
		14'b01000101001100: color_data = 12'b110011110111;
		14'b01000101001101: color_data = 12'b110011110111;
		14'b01000101001110: color_data = 12'b110011110111;
		14'b01000101010100: color_data = 12'b110011110111;
		14'b01000101010101: color_data = 12'b110011110111;
		14'b01000101010110: color_data = 12'b110011110111;
		14'b01000101010111: color_data = 12'b110011110111;
		14'b01000101011101: color_data = 12'b110011110111;
		14'b01000101011110: color_data = 12'b110011110111;
		14'b01000101011111: color_data = 12'b110011110111;
		14'b01000101100000: color_data = 12'b110011110111;
		14'b01000101100001: color_data = 12'b110011110111;
		14'b01000101101100: color_data = 12'b110011110111;
		14'b01000101101101: color_data = 12'b110011110111;
		14'b01000101101110: color_data = 12'b110011110111;
		14'b01000101101111: color_data = 12'b110011110111;
		14'b01000101110000: color_data = 12'b110011110111;
		14'b01000110000100: color_data = 12'b110011110111;
		14'b01000110000101: color_data = 12'b110011110111;
		14'b01000110000110: color_data = 12'b110011110111;
		14'b01000110000111: color_data = 12'b110011110111;
		14'b01000110001000: color_data = 12'b110011110111;
		14'b01000110001110: color_data = 12'b110011110111;
		14'b01000110001111: color_data = 12'b110011110111;
		14'b01000110010000: color_data = 12'b110011110111;
		14'b01000110010001: color_data = 12'b110011110111;
		14'b01000110010010: color_data = 12'b110011110111;
		14'b01000110011000: color_data = 12'b110011110111;
		14'b01000110011001: color_data = 12'b110011110111;
		14'b01000110011010: color_data = 12'b110011110111;
		14'b01000110011011: color_data = 12'b110011110111;
		14'b01000110011100: color_data = 12'b110011110111;
		14'b01000110100010: color_data = 12'b110011110111;
		14'b01000110100011: color_data = 12'b110011110111;
		14'b01000110100100: color_data = 12'b110011110111;
		14'b01000110100101: color_data = 12'b110011110111;
		14'b01000110100110: color_data = 12'b110011110111;
		14'b01000110101011: color_data = 12'b110011110111;
		14'b01000110101100: color_data = 12'b110011110111;
		14'b01000110101101: color_data = 12'b110011110111;
		14'b01000110101110: color_data = 12'b110011110111;
		14'b01000110101111: color_data = 12'b110011110111;
		14'b01000110110101: color_data = 12'b110011110111;
		14'b01000110110110: color_data = 12'b110011110111;
		14'b01000110110111: color_data = 12'b110011110111;
		14'b01000110111000: color_data = 12'b110011110111;
		14'b01000110111001: color_data = 12'b110011110111;
		14'b01000110111111: color_data = 12'b110011110111;
		14'b01000111000000: color_data = 12'b110011110111;
		14'b01000111000001: color_data = 12'b110011110111;
		14'b01000111000010: color_data = 12'b110011110111;
		14'b01000111000011: color_data = 12'b110011110111;
		14'b01000111001001: color_data = 12'b110011110111;
		14'b01000111001010: color_data = 12'b110011110111;
		14'b01000111001011: color_data = 12'b110011110111;
		14'b01000111001100: color_data = 12'b110011110111;
		14'b01000111001101: color_data = 12'b110011110111;
		14'b01001000001111: color_data = 12'b110011110111;
		14'b01001000010000: color_data = 12'b110011110111;
		14'b01001000010001: color_data = 12'b110011110111;
		14'b01001000010010: color_data = 12'b110011110111;
		14'b01001000010011: color_data = 12'b110011110111;
		14'b01001000011001: color_data = 12'b110011110111;
		14'b01001000011010: color_data = 12'b110011110111;
		14'b01001000011011: color_data = 12'b110011110111;
		14'b01001000011100: color_data = 12'b110011110111;
		14'b01001000011101: color_data = 12'b110011110111;
		14'b01001000100011: color_data = 12'b110011110111;
		14'b01001000100100: color_data = 12'b110011110111;
		14'b01001000100101: color_data = 12'b110011110111;
		14'b01001000100110: color_data = 12'b110011110111;
		14'b01001000100111: color_data = 12'b110011110111;
		14'b01001000101100: color_data = 12'b110011110111;
		14'b01001000101101: color_data = 12'b110011110111;
		14'b01001000101110: color_data = 12'b110011110111;
		14'b01001000101111: color_data = 12'b110011110111;
		14'b01001000110000: color_data = 12'b110011110111;
		14'b01001000110110: color_data = 12'b110011110111;
		14'b01001000110111: color_data = 12'b110011110111;
		14'b01001000111000: color_data = 12'b110011110111;
		14'b01001000111001: color_data = 12'b110011110111;
		14'b01001000111010: color_data = 12'b110011110111;
		14'b01001001000000: color_data = 12'b110011110111;
		14'b01001001000001: color_data = 12'b110011110111;
		14'b01001001000010: color_data = 12'b110011110111;
		14'b01001001000011: color_data = 12'b110011110111;
		14'b01001001000100: color_data = 12'b110011110111;
		14'b01001001001010: color_data = 12'b110011110111;
		14'b01001001001011: color_data = 12'b110011110111;
		14'b01001001001100: color_data = 12'b110011110111;
		14'b01001001001101: color_data = 12'b110011110111;
		14'b01001001001110: color_data = 12'b110011110111;
		14'b01001001010100: color_data = 12'b110011110111;
		14'b01001001010101: color_data = 12'b110011110111;
		14'b01001001010110: color_data = 12'b110011110111;
		14'b01001001010111: color_data = 12'b110011110111;
		14'b01001001011101: color_data = 12'b110011110111;
		14'b01001001011110: color_data = 12'b110011110111;
		14'b01001001011111: color_data = 12'b110011110111;
		14'b01001001100000: color_data = 12'b110011110111;
		14'b01001001100001: color_data = 12'b110011110111;
		14'b01001001101100: color_data = 12'b110011110111;
		14'b01001001101101: color_data = 12'b110011110111;
		14'b01001001101110: color_data = 12'b110011110111;
		14'b01001001101111: color_data = 12'b110011110111;
		14'b01001001110000: color_data = 12'b110011110111;
		14'b01001010000100: color_data = 12'b110011110111;
		14'b01001010000101: color_data = 12'b110011110111;
		14'b01001010000110: color_data = 12'b110011110111;
		14'b01001010000111: color_data = 12'b110011110111;
		14'b01001010001000: color_data = 12'b110011110111;
		14'b01001010001110: color_data = 12'b110011110111;
		14'b01001010001111: color_data = 12'b110011110111;
		14'b01001010010000: color_data = 12'b110011110111;
		14'b01001010010001: color_data = 12'b110011110111;
		14'b01001010010010: color_data = 12'b110011110111;
		14'b01001010011000: color_data = 12'b110011110111;
		14'b01001010011001: color_data = 12'b110011110111;
		14'b01001010011010: color_data = 12'b110011110111;
		14'b01001010011011: color_data = 12'b110011110111;
		14'b01001010011100: color_data = 12'b110011110111;
		14'b01001010100010: color_data = 12'b110011110111;
		14'b01001010100011: color_data = 12'b110011110111;
		14'b01001010100100: color_data = 12'b110011110111;
		14'b01001010100101: color_data = 12'b110011110111;
		14'b01001010100110: color_data = 12'b110011110111;
		14'b01001010101011: color_data = 12'b110011110111;
		14'b01001010101100: color_data = 12'b110011110111;
		14'b01001010101101: color_data = 12'b110011110111;
		14'b01001010101110: color_data = 12'b110011110111;
		14'b01001010101111: color_data = 12'b110011110111;
		14'b01001010110101: color_data = 12'b110011110111;
		14'b01001010110110: color_data = 12'b110011110111;
		14'b01001010110111: color_data = 12'b110011110111;
		14'b01001010111000: color_data = 12'b110011110111;
		14'b01001010111001: color_data = 12'b110011110111;
		14'b01001010111111: color_data = 12'b110011110111;
		14'b01001011000000: color_data = 12'b110011110111;
		14'b01001011000001: color_data = 12'b110011110111;
		14'b01001011000010: color_data = 12'b110011110111;
		14'b01001011000011: color_data = 12'b110011110111;
		14'b01001011001001: color_data = 12'b110011110111;
		14'b01001011001010: color_data = 12'b110011110111;
		14'b01001011001011: color_data = 12'b110011110111;
		14'b01001011001100: color_data = 12'b110011110111;
		14'b01001011001101: color_data = 12'b110011110111;
		14'b01001100000000: color_data = 12'b110011110111;
		14'b01001100000001: color_data = 12'b110011110111;
		14'b01001100000010: color_data = 12'b110011110111;
		14'b01001100000011: color_data = 12'b110011110111;
		14'b01001100000100: color_data = 12'b110011110111;
		14'b01001100000101: color_data = 12'b110011110111;
		14'b01001100000110: color_data = 12'b110011110111;
		14'b01001100000111: color_data = 12'b110011110111;
		14'b01001100001000: color_data = 12'b110011110111;
		14'b01001100001001: color_data = 12'b110011110111;
		14'b01001100001010: color_data = 12'b110011110111;
		14'b01001100001011: color_data = 12'b110011110111;
		14'b01001100001100: color_data = 12'b110011110111;
		14'b01001100001101: color_data = 12'b110011110111;
		14'b01001100001110: color_data = 12'b110011110111;
		14'b01001100001111: color_data = 12'b110011110111;
		14'b01001100010000: color_data = 12'b110011110111;
		14'b01001100010001: color_data = 12'b110011110111;
		14'b01001100010010: color_data = 12'b110011110111;
		14'b01001100010011: color_data = 12'b110011110111;
		14'b01001100011001: color_data = 12'b110011110111;
		14'b01001100011010: color_data = 12'b110011110111;
		14'b01001100011011: color_data = 12'b110011110111;
		14'b01001100011100: color_data = 12'b110011110111;
		14'b01001100011101: color_data = 12'b110011110111;
		14'b01001100100011: color_data = 12'b110011110111;
		14'b01001100100100: color_data = 12'b110011110111;
		14'b01001100100101: color_data = 12'b110011110111;
		14'b01001100100110: color_data = 12'b110011110111;
		14'b01001100100111: color_data = 12'b110011110111;
		14'b01001100101100: color_data = 12'b110011110111;
		14'b01001100101101: color_data = 12'b110011110111;
		14'b01001100101110: color_data = 12'b110011110111;
		14'b01001100101111: color_data = 12'b110011110111;
		14'b01001100110000: color_data = 12'b110011110111;
		14'b01001100110110: color_data = 12'b110011110111;
		14'b01001100110111: color_data = 12'b110011110111;
		14'b01001100111000: color_data = 12'b110011110111;
		14'b01001100111001: color_data = 12'b110011110111;
		14'b01001100111010: color_data = 12'b110011110111;
		14'b01001100111011: color_data = 12'b110011110111;
		14'b01001100111100: color_data = 12'b110011110111;
		14'b01001100111101: color_data = 12'b110011110111;
		14'b01001100111110: color_data = 12'b110011110111;
		14'b01001100111111: color_data = 12'b110011110111;
		14'b01001101000000: color_data = 12'b110011110111;
		14'b01001101000001: color_data = 12'b110011110111;
		14'b01001101000010: color_data = 12'b110011110111;
		14'b01001101000011: color_data = 12'b110011110111;
		14'b01001101000100: color_data = 12'b110011110111;
		14'b01001101001010: color_data = 12'b110011110111;
		14'b01001101001011: color_data = 12'b110011110111;
		14'b01001101001100: color_data = 12'b110011110111;
		14'b01001101001101: color_data = 12'b110011110111;
		14'b01001101001110: color_data = 12'b110011110111;
		14'b01001101010100: color_data = 12'b110011110111;
		14'b01001101010101: color_data = 12'b110011110111;
		14'b01001101010110: color_data = 12'b110011110111;
		14'b01001101010111: color_data = 12'b110011110111;
		14'b01001101011000: color_data = 12'b110011110111;
		14'b01001101011001: color_data = 12'b110011110111;
		14'b01001101011010: color_data = 12'b110011110111;
		14'b01001101011011: color_data = 12'b110011110111;
		14'b01001101011100: color_data = 12'b110011110111;
		14'b01001101101100: color_data = 12'b110011110111;
		14'b01001101101101: color_data = 12'b110011110111;
		14'b01001101101110: color_data = 12'b110011110111;
		14'b01001101101111: color_data = 12'b110011110111;
		14'b01001101110000: color_data = 12'b110011110111;
		14'b01001110000100: color_data = 12'b110011110111;
		14'b01001110000101: color_data = 12'b110011110111;
		14'b01001110000110: color_data = 12'b110011110111;
		14'b01001110000111: color_data = 12'b110011110111;
		14'b01001110001000: color_data = 12'b110011110111;
		14'b01001110001110: color_data = 12'b110011110111;
		14'b01001110001111: color_data = 12'b110011110111;
		14'b01001110010000: color_data = 12'b110011110111;
		14'b01001110010001: color_data = 12'b110011110111;
		14'b01001110010010: color_data = 12'b110011110111;
		14'b01001110010011: color_data = 12'b110011110111;
		14'b01001110010100: color_data = 12'b110011110111;
		14'b01001110010101: color_data = 12'b110011110111;
		14'b01001110010110: color_data = 12'b110011110111;
		14'b01001110010111: color_data = 12'b110011110111;
		14'b01001110011000: color_data = 12'b110011110111;
		14'b01001110011001: color_data = 12'b110011110111;
		14'b01001110011010: color_data = 12'b110011110111;
		14'b01001110011011: color_data = 12'b110011110111;
		14'b01001110011100: color_data = 12'b110011110111;
		14'b01001110100010: color_data = 12'b110011110111;
		14'b01001110100011: color_data = 12'b110011110111;
		14'b01001110100100: color_data = 12'b110011110111;
		14'b01001110100101: color_data = 12'b110011110111;
		14'b01001110100110: color_data = 12'b110011110111;
		14'b01001110100111: color_data = 12'b110011110111;
		14'b01001110101000: color_data = 12'b110011110111;
		14'b01001110101001: color_data = 12'b110011110111;
		14'b01001110101010: color_data = 12'b110011110111;
		14'b01001110101011: color_data = 12'b110011110111;
		14'b01001110101100: color_data = 12'b110011110111;
		14'b01001110101101: color_data = 12'b110011110111;
		14'b01001110101110: color_data = 12'b110011110111;
		14'b01001110101111: color_data = 12'b110011110111;
		14'b01001110110101: color_data = 12'b110011110111;
		14'b01001110110110: color_data = 12'b110011110111;
		14'b01001110110111: color_data = 12'b110011110111;
		14'b01001110111000: color_data = 12'b110011110111;
		14'b01001110111001: color_data = 12'b110011110111;
		14'b01001110111010: color_data = 12'b110011110111;
		14'b01001110111011: color_data = 12'b110011110111;
		14'b01001110111100: color_data = 12'b110011110111;
		14'b01001110111101: color_data = 12'b110011110111;
		14'b01001110111110: color_data = 12'b110011110111;
		14'b01001111001001: color_data = 12'b110011110111;
		14'b01001111001010: color_data = 12'b110011110111;
		14'b01001111001011: color_data = 12'b110011110111;
		14'b01001111001100: color_data = 12'b110011110111;
		14'b01001111001101: color_data = 12'b110011110111;
		14'b01010000000000: color_data = 12'b110011110111;
		14'b01010000000001: color_data = 12'b110011110111;
		14'b01010000000010: color_data = 12'b110011110111;
		14'b01010000000011: color_data = 12'b110011110111;
		14'b01010000000100: color_data = 12'b110011110111;
		14'b01010000000101: color_data = 12'b110011110111;
		14'b01010000000110: color_data = 12'b110011110111;
		14'b01010000000111: color_data = 12'b110011110111;
		14'b01010000001000: color_data = 12'b110011110111;
		14'b01010000001001: color_data = 12'b110011110111;
		14'b01010000001010: color_data = 12'b110011110111;
		14'b01010000001011: color_data = 12'b110011110111;
		14'b01010000001100: color_data = 12'b110011110111;
		14'b01010000001101: color_data = 12'b110011110111;
		14'b01010000001110: color_data = 12'b110011110111;
		14'b01010000001111: color_data = 12'b110011110111;
		14'b01010000010000: color_data = 12'b110011110111;
		14'b01010000010001: color_data = 12'b110011110111;
		14'b01010000010010: color_data = 12'b110011110111;
		14'b01010000010011: color_data = 12'b110011110111;
		14'b01010000011001: color_data = 12'b110011110111;
		14'b01010000011010: color_data = 12'b110011110111;
		14'b01010000011011: color_data = 12'b110011110111;
		14'b01010000011100: color_data = 12'b110011110111;
		14'b01010000011101: color_data = 12'b110011110111;
		14'b01010000100011: color_data = 12'b110011110111;
		14'b01010000100100: color_data = 12'b110011110111;
		14'b01010000100101: color_data = 12'b110011110111;
		14'b01010000100110: color_data = 12'b110011110111;
		14'b01010000100111: color_data = 12'b110011110111;
		14'b01010000101100: color_data = 12'b110011110111;
		14'b01010000101101: color_data = 12'b110011110111;
		14'b01010000101110: color_data = 12'b110011110111;
		14'b01010000101111: color_data = 12'b110011110111;
		14'b01010000110000: color_data = 12'b110011110111;
		14'b01010000110110: color_data = 12'b110011110111;
		14'b01010000110111: color_data = 12'b110011110111;
		14'b01010000111000: color_data = 12'b110011110111;
		14'b01010000111001: color_data = 12'b110011110111;
		14'b01010000111010: color_data = 12'b110011110111;
		14'b01010000111011: color_data = 12'b110011110111;
		14'b01010000111100: color_data = 12'b110011110111;
		14'b01010000111101: color_data = 12'b110011110111;
		14'b01010000111110: color_data = 12'b110011110111;
		14'b01010000111111: color_data = 12'b110011110111;
		14'b01010001000000: color_data = 12'b110011110111;
		14'b01010001000001: color_data = 12'b110011110111;
		14'b01010001000010: color_data = 12'b110011110111;
		14'b01010001000011: color_data = 12'b110011110111;
		14'b01010001000100: color_data = 12'b110011110111;
		14'b01010001001010: color_data = 12'b110011110111;
		14'b01010001001011: color_data = 12'b110011110111;
		14'b01010001001100: color_data = 12'b110011110111;
		14'b01010001001101: color_data = 12'b110011110111;
		14'b01010001001110: color_data = 12'b110011110111;
		14'b01010001010100: color_data = 12'b110011110111;
		14'b01010001010101: color_data = 12'b110011110111;
		14'b01010001010110: color_data = 12'b110011110111;
		14'b01010001010111: color_data = 12'b110011110111;
		14'b01010001011000: color_data = 12'b110011110111;
		14'b01010001011001: color_data = 12'b110011110111;
		14'b01010001011010: color_data = 12'b110011110111;
		14'b01010001011011: color_data = 12'b110011110111;
		14'b01010001011100: color_data = 12'b110011110111;
		14'b01010001101100: color_data = 12'b110011110111;
		14'b01010001101101: color_data = 12'b110011110111;
		14'b01010001101110: color_data = 12'b110011110111;
		14'b01010001101111: color_data = 12'b110011110111;
		14'b01010001110000: color_data = 12'b110011110111;
		14'b01010010000100: color_data = 12'b110011110111;
		14'b01010010000101: color_data = 12'b110011110111;
		14'b01010010000110: color_data = 12'b110011110111;
		14'b01010010000111: color_data = 12'b110011110111;
		14'b01010010001000: color_data = 12'b110011110111;
		14'b01010010001110: color_data = 12'b110011110111;
		14'b01010010001111: color_data = 12'b110011110111;
		14'b01010010010000: color_data = 12'b110011110111;
		14'b01010010010001: color_data = 12'b110011110111;
		14'b01010010010010: color_data = 12'b110011110111;
		14'b01010010010011: color_data = 12'b110011110111;
		14'b01010010010100: color_data = 12'b110011110111;
		14'b01010010010101: color_data = 12'b110011110111;
		14'b01010010010110: color_data = 12'b110011110111;
		14'b01010010010111: color_data = 12'b110011110111;
		14'b01010010011000: color_data = 12'b110011110111;
		14'b01010010011001: color_data = 12'b110011110111;
		14'b01010010011010: color_data = 12'b110011110111;
		14'b01010010011011: color_data = 12'b110011110111;
		14'b01010010011100: color_data = 12'b110011110111;
		14'b01010010100010: color_data = 12'b110011110111;
		14'b01010010100011: color_data = 12'b110011110111;
		14'b01010010100100: color_data = 12'b110011110111;
		14'b01010010100101: color_data = 12'b110011110111;
		14'b01010010100110: color_data = 12'b110011110111;
		14'b01010010100111: color_data = 12'b110011110111;
		14'b01010010101000: color_data = 12'b110011110111;
		14'b01010010101001: color_data = 12'b110011110111;
		14'b01010010101010: color_data = 12'b110011110111;
		14'b01010010101011: color_data = 12'b110011110111;
		14'b01010010101100: color_data = 12'b110011110111;
		14'b01010010101101: color_data = 12'b110011110111;
		14'b01010010101110: color_data = 12'b110011110111;
		14'b01010010101111: color_data = 12'b110011110111;
		14'b01010010110101: color_data = 12'b110011110111;
		14'b01010010110110: color_data = 12'b110011110111;
		14'b01010010110111: color_data = 12'b110011110111;
		14'b01010010111000: color_data = 12'b110011110111;
		14'b01010010111001: color_data = 12'b110011110111;
		14'b01010010111010: color_data = 12'b110011110111;
		14'b01010010111011: color_data = 12'b110011110111;
		14'b01010010111100: color_data = 12'b110011110111;
		14'b01010010111101: color_data = 12'b110011110111;
		14'b01010010111110: color_data = 12'b110011110111;
		14'b01010011001001: color_data = 12'b110011110111;
		14'b01010011001010: color_data = 12'b110011110111;
		14'b01010011001011: color_data = 12'b110011110111;
		14'b01010011001100: color_data = 12'b110011110111;
		14'b01010011001101: color_data = 12'b110011110111;
		14'b01010100000000: color_data = 12'b110011110111;
		14'b01010100000001: color_data = 12'b110011110111;
		14'b01010100000010: color_data = 12'b110011110111;
		14'b01010100000011: color_data = 12'b110011110111;
		14'b01010100000100: color_data = 12'b110011110111;
		14'b01010100000101: color_data = 12'b110011110111;
		14'b01010100000110: color_data = 12'b110011110111;
		14'b01010100000111: color_data = 12'b110011110111;
		14'b01010100001000: color_data = 12'b110011110111;
		14'b01010100001001: color_data = 12'b110011110111;
		14'b01010100001010: color_data = 12'b110011110111;
		14'b01010100001011: color_data = 12'b110011110111;
		14'b01010100001100: color_data = 12'b110011110111;
		14'b01010100001101: color_data = 12'b110011110111;
		14'b01010100001110: color_data = 12'b110011110111;
		14'b01010100001111: color_data = 12'b110011110111;
		14'b01010100010000: color_data = 12'b110011110111;
		14'b01010100010001: color_data = 12'b110011110111;
		14'b01010100010010: color_data = 12'b110011110111;
		14'b01010100010011: color_data = 12'b110011110111;
		14'b01010100011001: color_data = 12'b110011110111;
		14'b01010100011010: color_data = 12'b110011110111;
		14'b01010100011011: color_data = 12'b110011110111;
		14'b01010100011100: color_data = 12'b110011110111;
		14'b01010100011101: color_data = 12'b110011110111;
		14'b01010100100011: color_data = 12'b110011110111;
		14'b01010100100100: color_data = 12'b110011110111;
		14'b01010100100101: color_data = 12'b110011110111;
		14'b01010100100110: color_data = 12'b110011110111;
		14'b01010100100111: color_data = 12'b110011110111;
		14'b01010100101100: color_data = 12'b110011110111;
		14'b01010100101101: color_data = 12'b110011110111;
		14'b01010100101110: color_data = 12'b110011110111;
		14'b01010100101111: color_data = 12'b110011110111;
		14'b01010100110000: color_data = 12'b110011110111;
		14'b01010100110110: color_data = 12'b110011110111;
		14'b01010100110111: color_data = 12'b110011110111;
		14'b01010100111000: color_data = 12'b110011110111;
		14'b01010100111001: color_data = 12'b110011110111;
		14'b01010100111010: color_data = 12'b110011110111;
		14'b01010100111011: color_data = 12'b110011110111;
		14'b01010100111100: color_data = 12'b110011110111;
		14'b01010100111101: color_data = 12'b110011110111;
		14'b01010100111110: color_data = 12'b110011110111;
		14'b01010100111111: color_data = 12'b110011110111;
		14'b01010101000000: color_data = 12'b110011110111;
		14'b01010101000001: color_data = 12'b110011110111;
		14'b01010101000010: color_data = 12'b110011110111;
		14'b01010101000011: color_data = 12'b110011110111;
		14'b01010101000100: color_data = 12'b110011110111;
		14'b01010101001010: color_data = 12'b110011110111;
		14'b01010101001011: color_data = 12'b110011110111;
		14'b01010101001100: color_data = 12'b110011110111;
		14'b01010101001101: color_data = 12'b110011110111;
		14'b01010101001110: color_data = 12'b110011110111;
		14'b01010101010100: color_data = 12'b110011110111;
		14'b01010101010101: color_data = 12'b110011110111;
		14'b01010101010110: color_data = 12'b110011110111;
		14'b01010101010111: color_data = 12'b110011110111;
		14'b01010101011000: color_data = 12'b110011110111;
		14'b01010101011001: color_data = 12'b110011110111;
		14'b01010101011010: color_data = 12'b110011110111;
		14'b01010101011011: color_data = 12'b110011110111;
		14'b01010101011100: color_data = 12'b110011110111;
		14'b01010101101100: color_data = 12'b110011110111;
		14'b01010101101101: color_data = 12'b110011110111;
		14'b01010101101110: color_data = 12'b110011110111;
		14'b01010101101111: color_data = 12'b110011110111;
		14'b01010101110000: color_data = 12'b110011110111;
		14'b01010110000100: color_data = 12'b110011110111;
		14'b01010110000101: color_data = 12'b110011110111;
		14'b01010110000110: color_data = 12'b110011110111;
		14'b01010110000111: color_data = 12'b110011110111;
		14'b01010110001000: color_data = 12'b110011110111;
		14'b01010110001110: color_data = 12'b110011110111;
		14'b01010110001111: color_data = 12'b110011110111;
		14'b01010110010000: color_data = 12'b110011110111;
		14'b01010110010001: color_data = 12'b110011110111;
		14'b01010110010010: color_data = 12'b110011110111;
		14'b01010110010011: color_data = 12'b110011110111;
		14'b01010110010100: color_data = 12'b110011110111;
		14'b01010110010101: color_data = 12'b110011110111;
		14'b01010110010110: color_data = 12'b110011110111;
		14'b01010110010111: color_data = 12'b110011110111;
		14'b01010110011000: color_data = 12'b110011110111;
		14'b01010110011001: color_data = 12'b110011110111;
		14'b01010110011010: color_data = 12'b110011110111;
		14'b01010110011011: color_data = 12'b110011110111;
		14'b01010110011100: color_data = 12'b110011110111;
		14'b01010110100010: color_data = 12'b110011110111;
		14'b01010110100011: color_data = 12'b110011110111;
		14'b01010110100100: color_data = 12'b110011110111;
		14'b01010110100101: color_data = 12'b110011110111;
		14'b01010110100110: color_data = 12'b110011110111;
		14'b01010110100111: color_data = 12'b110011110111;
		14'b01010110101000: color_data = 12'b110011110111;
		14'b01010110101001: color_data = 12'b110011110111;
		14'b01010110101010: color_data = 12'b110011110111;
		14'b01010110101011: color_data = 12'b110011110111;
		14'b01010110101100: color_data = 12'b110011110111;
		14'b01010110101101: color_data = 12'b110011110111;
		14'b01010110101110: color_data = 12'b110011110111;
		14'b01010110101111: color_data = 12'b110011110111;
		14'b01010110110101: color_data = 12'b110011110111;
		14'b01010110110110: color_data = 12'b110011110111;
		14'b01010110110111: color_data = 12'b110011110111;
		14'b01010110111000: color_data = 12'b110011110111;
		14'b01010110111001: color_data = 12'b110011110111;
		14'b01010110111010: color_data = 12'b110011110111;
		14'b01010110111011: color_data = 12'b110011110111;
		14'b01010110111100: color_data = 12'b110011110111;
		14'b01010110111101: color_data = 12'b110011110111;
		14'b01010110111110: color_data = 12'b110011110111;
		14'b01010111001001: color_data = 12'b110011110111;
		14'b01010111001010: color_data = 12'b110011110111;
		14'b01010111001011: color_data = 12'b110011110111;
		14'b01010111001100: color_data = 12'b110011110111;
		14'b01010111001101: color_data = 12'b110011110111;
		14'b01011000000000: color_data = 12'b110011110111;
		14'b01011000000001: color_data = 12'b110011110111;
		14'b01011000000010: color_data = 12'b110011110111;
		14'b01011000000011: color_data = 12'b110011110111;
		14'b01011000000100: color_data = 12'b110011110111;
		14'b01011000000101: color_data = 12'b110011110111;
		14'b01011000000110: color_data = 12'b110011110111;
		14'b01011000000111: color_data = 12'b110011110111;
		14'b01011000001000: color_data = 12'b110011110111;
		14'b01011000001001: color_data = 12'b110011110111;
		14'b01011000001010: color_data = 12'b110011110111;
		14'b01011000001011: color_data = 12'b110011110111;
		14'b01011000001100: color_data = 12'b110011110111;
		14'b01011000001101: color_data = 12'b110011110111;
		14'b01011000001110: color_data = 12'b110011110111;
		14'b01011000001111: color_data = 12'b110011110111;
		14'b01011000010000: color_data = 12'b110011110111;
		14'b01011000010001: color_data = 12'b110011110111;
		14'b01011000010010: color_data = 12'b110011110111;
		14'b01011000010011: color_data = 12'b110011110111;
		14'b01011000011001: color_data = 12'b110011110111;
		14'b01011000011010: color_data = 12'b110011110111;
		14'b01011000011011: color_data = 12'b110011110111;
		14'b01011000011100: color_data = 12'b110011110111;
		14'b01011000011101: color_data = 12'b110011110111;
		14'b01011000100011: color_data = 12'b110011110111;
		14'b01011000100100: color_data = 12'b110011110111;
		14'b01011000100101: color_data = 12'b110011110111;
		14'b01011000100110: color_data = 12'b110011110111;
		14'b01011000100111: color_data = 12'b110011110111;
		14'b01011000101100: color_data = 12'b110011110111;
		14'b01011000101101: color_data = 12'b110011110111;
		14'b01011000101110: color_data = 12'b110011110111;
		14'b01011000101111: color_data = 12'b110011110111;
		14'b01011000110000: color_data = 12'b110011110111;
		14'b01011000110110: color_data = 12'b110011110111;
		14'b01011000110111: color_data = 12'b110011110111;
		14'b01011000111000: color_data = 12'b110011110111;
		14'b01011000111001: color_data = 12'b110011110111;
		14'b01011000111010: color_data = 12'b110011110111;
		14'b01011000111011: color_data = 12'b110011110111;
		14'b01011000111100: color_data = 12'b110011110111;
		14'b01011000111101: color_data = 12'b110011110111;
		14'b01011000111110: color_data = 12'b110011110111;
		14'b01011000111111: color_data = 12'b110011110111;
		14'b01011001000000: color_data = 12'b110011110111;
		14'b01011001000001: color_data = 12'b110011110111;
		14'b01011001000010: color_data = 12'b110011110111;
		14'b01011001000011: color_data = 12'b110011110111;
		14'b01011001000100: color_data = 12'b110011110111;
		14'b01011001001010: color_data = 12'b110011110111;
		14'b01011001001011: color_data = 12'b110011110111;
		14'b01011001001100: color_data = 12'b110011110111;
		14'b01011001001101: color_data = 12'b110011110111;
		14'b01011001001110: color_data = 12'b110011110111;
		14'b01011001010100: color_data = 12'b110011110111;
		14'b01011001010101: color_data = 12'b110011110111;
		14'b01011001010110: color_data = 12'b110011110111;
		14'b01011001010111: color_data = 12'b110011110111;
		14'b01011001011000: color_data = 12'b110011110111;
		14'b01011001011001: color_data = 12'b110011110111;
		14'b01011001011010: color_data = 12'b110011110111;
		14'b01011001011011: color_data = 12'b110011110111;
		14'b01011001011100: color_data = 12'b110011110111;
		14'b01011001101100: color_data = 12'b110011110111;
		14'b01011001101101: color_data = 12'b110011110111;
		14'b01011001101110: color_data = 12'b110011110111;
		14'b01011001101111: color_data = 12'b110011110111;
		14'b01011001110000: color_data = 12'b110011110111;
		14'b01011010000100: color_data = 12'b110011110111;
		14'b01011010000101: color_data = 12'b110011110111;
		14'b01011010000110: color_data = 12'b110011110111;
		14'b01011010000111: color_data = 12'b110011110111;
		14'b01011010001000: color_data = 12'b110011110111;
		14'b01011010001110: color_data = 12'b110011110111;
		14'b01011010001111: color_data = 12'b110011110111;
		14'b01011010010000: color_data = 12'b110011110111;
		14'b01011010010001: color_data = 12'b110011110111;
		14'b01011010010010: color_data = 12'b110011110111;
		14'b01011010010011: color_data = 12'b110011110111;
		14'b01011010010100: color_data = 12'b110011110111;
		14'b01011010010101: color_data = 12'b110011110111;
		14'b01011010010110: color_data = 12'b110011110111;
		14'b01011010010111: color_data = 12'b110011110111;
		14'b01011010011000: color_data = 12'b110011110111;
		14'b01011010011001: color_data = 12'b110011110111;
		14'b01011010011010: color_data = 12'b110011110111;
		14'b01011010011011: color_data = 12'b110011110111;
		14'b01011010011100: color_data = 12'b110011110111;
		14'b01011010100010: color_data = 12'b110011110111;
		14'b01011010100011: color_data = 12'b110011110111;
		14'b01011010100100: color_data = 12'b110011110111;
		14'b01011010100101: color_data = 12'b110011110111;
		14'b01011010100110: color_data = 12'b110011110111;
		14'b01011010100111: color_data = 12'b110011110111;
		14'b01011010101000: color_data = 12'b110011110111;
		14'b01011010101001: color_data = 12'b110011110111;
		14'b01011010101010: color_data = 12'b110011110111;
		14'b01011010101011: color_data = 12'b110011110111;
		14'b01011010101100: color_data = 12'b110011110111;
		14'b01011010101101: color_data = 12'b110011110111;
		14'b01011010101110: color_data = 12'b110011110111;
		14'b01011010101111: color_data = 12'b110011110111;
		14'b01011010110101: color_data = 12'b110011110111;
		14'b01011010110110: color_data = 12'b110011110111;
		14'b01011010110111: color_data = 12'b110011110111;
		14'b01011010111000: color_data = 12'b110011110111;
		14'b01011010111001: color_data = 12'b110011110111;
		14'b01011010111010: color_data = 12'b110011110111;
		14'b01011010111011: color_data = 12'b110011110111;
		14'b01011010111100: color_data = 12'b110011110111;
		14'b01011010111101: color_data = 12'b110011110111;
		14'b01011010111110: color_data = 12'b110011110111;
		14'b01011011001001: color_data = 12'b110011110111;
		14'b01011011001010: color_data = 12'b110011110111;
		14'b01011011001011: color_data = 12'b110011110111;
		14'b01011011001100: color_data = 12'b110011110111;
		14'b01011011001101: color_data = 12'b110011110111;
		14'b01011101000000: color_data = 12'b110011110111;
		14'b01011101000001: color_data = 12'b110011110111;
		14'b01011101000010: color_data = 12'b110011110111;
		14'b01011101000011: color_data = 12'b110011110111;
		14'b01011101000100: color_data = 12'b110011110111;
		14'b01011110101011: color_data = 12'b110011110111;
		14'b01011110101100: color_data = 12'b110011110111;
		14'b01011110101101: color_data = 12'b110011110111;
		14'b01011110101110: color_data = 12'b110011110111;
		14'b01011110101111: color_data = 12'b110011110111;
		14'b01100001000000: color_data = 12'b110011110111;
		14'b01100001000001: color_data = 12'b110011110111;
		14'b01100001000010: color_data = 12'b110011110111;
		14'b01100001000011: color_data = 12'b110011110111;
		14'b01100001000100: color_data = 12'b110011110111;
		14'b01100010101011: color_data = 12'b110011110111;
		14'b01100010101100: color_data = 12'b110011110111;
		14'b01100010101101: color_data = 12'b110011110111;
		14'b01100010101110: color_data = 12'b110011110111;
		14'b01100010101111: color_data = 12'b110011110111;
		14'b01100101000000: color_data = 12'b110011110111;
		14'b01100101000001: color_data = 12'b110011110111;
		14'b01100101000010: color_data = 12'b110011110111;
		14'b01100101000011: color_data = 12'b110011110111;
		14'b01100101000100: color_data = 12'b110011110111;
		14'b01100110101011: color_data = 12'b110011110111;
		14'b01100110101100: color_data = 12'b110011110111;
		14'b01100110101101: color_data = 12'b110011110111;
		14'b01100110101110: color_data = 12'b110011110111;
		14'b01100110101111: color_data = 12'b110011110111;
		14'b01101001000000: color_data = 12'b110011110111;
		14'b01101001000001: color_data = 12'b110011110111;
		14'b01101001000010: color_data = 12'b110011110111;
		14'b01101001000011: color_data = 12'b110011110111;
		14'b01101001000100: color_data = 12'b110011110111;
		14'b01101010101011: color_data = 12'b110011110111;
		14'b01101010101100: color_data = 12'b110011110111;
		14'b01101010101101: color_data = 12'b110011110111;
		14'b01101010101110: color_data = 12'b110011110111;
		14'b01101010101111: color_data = 12'b110011110111;
		14'b01101101000000: color_data = 12'b110011110111;
		14'b01101101000001: color_data = 12'b110011110111;
		14'b01101101000010: color_data = 12'b110011110111;
		14'b01101101000011: color_data = 12'b110011110111;
		14'b01101101000100: color_data = 12'b110011110111;
		14'b01101110101011: color_data = 12'b110011110111;
		14'b01101110101100: color_data = 12'b110011110111;
		14'b01101110101101: color_data = 12'b110011110111;
		14'b01101110101110: color_data = 12'b110011110111;
		14'b01101110101111: color_data = 12'b110011110111;
		14'b01110000110110: color_data = 12'b110011110111;
		14'b01110000110111: color_data = 12'b110011110111;
		14'b01110000111000: color_data = 12'b110011110111;
		14'b01110000111001: color_data = 12'b110011110111;
		14'b01110000111010: color_data = 12'b110011110111;
		14'b01110000111011: color_data = 12'b110011110111;
		14'b01110000111100: color_data = 12'b110011110111;
		14'b01110000111101: color_data = 12'b110011110111;
		14'b01110000111110: color_data = 12'b110011110111;
		14'b01110000111111: color_data = 12'b110011110111;
		14'b01110001000000: color_data = 12'b110011110111;
		14'b01110001000001: color_data = 12'b110011110111;
		14'b01110001000010: color_data = 12'b110011110111;
		14'b01110001000011: color_data = 12'b110011110111;
		14'b01110001000100: color_data = 12'b110011110111;
		14'b01110010100010: color_data = 12'b110011110111;
		14'b01110010100011: color_data = 12'b110011110111;
		14'b01110010100100: color_data = 12'b110011110111;
		14'b01110010100101: color_data = 12'b110011110111;
		14'b01110010100110: color_data = 12'b110011110111;
		14'b01110010100111: color_data = 12'b110011110111;
		14'b01110010101000: color_data = 12'b110011110111;
		14'b01110010101001: color_data = 12'b110011110111;
		14'b01110010101010: color_data = 12'b110011110111;
		14'b01110010101011: color_data = 12'b110011110111;
		14'b01110010101100: color_data = 12'b110011110111;
		14'b01110010101101: color_data = 12'b110011110111;
		14'b01110010101110: color_data = 12'b110011110111;
		14'b01110010101111: color_data = 12'b110011110111;
		14'b01110100110110: color_data = 12'b110011110111;
		14'b01110100110111: color_data = 12'b110011110111;
		14'b01110100111000: color_data = 12'b110011110111;
		14'b01110100111001: color_data = 12'b110011110111;
		14'b01110100111010: color_data = 12'b110011110111;
		14'b01110100111011: color_data = 12'b110011110111;
		14'b01110100111100: color_data = 12'b110011110111;
		14'b01110100111101: color_data = 12'b110011110111;
		14'b01110100111110: color_data = 12'b110011110111;
		14'b01110100111111: color_data = 12'b110011110111;
		14'b01110101000000: color_data = 12'b110011110111;
		14'b01110101000001: color_data = 12'b110011110111;
		14'b01110101000010: color_data = 12'b110011110111;
		14'b01110101000011: color_data = 12'b110011110111;
		14'b01110101000100: color_data = 12'b110011110111;
		14'b01110110100010: color_data = 12'b110011110111;
		14'b01110110100011: color_data = 12'b110011110111;
		14'b01110110100100: color_data = 12'b110011110111;
		14'b01110110100101: color_data = 12'b110011110111;
		14'b01110110100110: color_data = 12'b110011110111;
		14'b01110110100111: color_data = 12'b110011110111;
		14'b01110110101000: color_data = 12'b110011110111;
		14'b01110110101001: color_data = 12'b110011110111;
		14'b01110110101010: color_data = 12'b110011110111;
		14'b01110110101011: color_data = 12'b110011110111;
		14'b01110110101100: color_data = 12'b110011110111;
		14'b01110110101101: color_data = 12'b110011110111;
		14'b01110110101110: color_data = 12'b110011110111;
		14'b01110110101111: color_data = 12'b110011110111;
		14'b01111000110110: color_data = 12'b110011110111;
		14'b01111000110111: color_data = 12'b110011110111;
		14'b01111000111000: color_data = 12'b110011110111;
		14'b01111000111001: color_data = 12'b110011110111;
		14'b01111000111010: color_data = 12'b110011110111;
		14'b01111000111011: color_data = 12'b110011110111;
		14'b01111000111100: color_data = 12'b110011110111;
		14'b01111000111101: color_data = 12'b110011110111;
		14'b01111000111110: color_data = 12'b110011110111;
		14'b01111000111111: color_data = 12'b110011110111;
		14'b01111001000000: color_data = 12'b110011110111;
		14'b01111001000001: color_data = 12'b110011110111;
		14'b01111001000010: color_data = 12'b110011110111;
		14'b01111001000011: color_data = 12'b110011110111;
		14'b01111001000100: color_data = 12'b110011110111;
		14'b01111010100010: color_data = 12'b110011110111;
		14'b01111010100011: color_data = 12'b110011110111;
		14'b01111010100100: color_data = 12'b110011110111;
		14'b01111010100101: color_data = 12'b110011110111;
		14'b01111010100110: color_data = 12'b110011110111;
		14'b01111010100111: color_data = 12'b110011110111;
		14'b01111010101000: color_data = 12'b110011110111;
		14'b01111010101001: color_data = 12'b110011110111;
		14'b01111010101010: color_data = 12'b110011110111;
		14'b01111010101011: color_data = 12'b110011110111;
		14'b01111010101100: color_data = 12'b110011110111;
		14'b01111010101101: color_data = 12'b110011110111;
		14'b01111010101110: color_data = 12'b110011110111;
		14'b01111010101111: color_data = 12'b110011110111;
		14'b01111100110110: color_data = 12'b110011110111;
		14'b01111100110111: color_data = 12'b110011110111;
		14'b01111100111000: color_data = 12'b110011110111;
		14'b01111100111001: color_data = 12'b110011110111;
		14'b01111100111010: color_data = 12'b110011110111;
		14'b01111100111011: color_data = 12'b110011110111;
		14'b01111100111100: color_data = 12'b110011110111;
		14'b01111100111101: color_data = 12'b110011110111;
		14'b01111100111110: color_data = 12'b110011110111;
		14'b01111100111111: color_data = 12'b110011110111;
		14'b01111101000000: color_data = 12'b110011110111;
		14'b01111101000001: color_data = 12'b110011110111;
		14'b01111101000010: color_data = 12'b110011110111;
		14'b01111101000011: color_data = 12'b110011110111;
		14'b01111101000100: color_data = 12'b110011110111;
		14'b01111110100010: color_data = 12'b110011110111;
		14'b01111110100011: color_data = 12'b110011110111;
		14'b01111110100100: color_data = 12'b110011110111;
		14'b01111110100101: color_data = 12'b110011110111;
		14'b01111110100110: color_data = 12'b110011110111;
		14'b01111110100111: color_data = 12'b110011110111;
		14'b01111110101000: color_data = 12'b110011110111;
		14'b01111110101001: color_data = 12'b110011110111;
		14'b01111110101010: color_data = 12'b110011110111;
		14'b01111110101011: color_data = 12'b110011110111;
		14'b01111110101100: color_data = 12'b110011110111;
		14'b01111110101101: color_data = 12'b110011110111;
		14'b01111110101110: color_data = 12'b110011110111;
		14'b01111110101111: color_data = 12'b110011110111;
		14'b10000000110110: color_data = 12'b110011110111;
		14'b10000000110111: color_data = 12'b110011110111;
		14'b10000000111000: color_data = 12'b110011110111;
		14'b10000000111001: color_data = 12'b110011110111;
		14'b10000000111010: color_data = 12'b110011110111;
		14'b10000000111011: color_data = 12'b110011110111;
		14'b10000000111100: color_data = 12'b110011110111;
		14'b10000000111101: color_data = 12'b110011110111;
		14'b10000000111110: color_data = 12'b110011110111;
		14'b10000000111111: color_data = 12'b110011110111;
		14'b10000001000000: color_data = 12'b110011110111;
		14'b10000001000001: color_data = 12'b110011110111;
		14'b10000001000010: color_data = 12'b110011110111;
		14'b10000001000011: color_data = 12'b110011110111;
		14'b10000001000100: color_data = 12'b110011110111;
		14'b10000010100010: color_data = 12'b110011110111;
		14'b10000010100011: color_data = 12'b110011110111;
		14'b10000010100100: color_data = 12'b110011110111;
		14'b10000010100101: color_data = 12'b110011110111;
		14'b10000010100110: color_data = 12'b110011110111;
		14'b10000010100111: color_data = 12'b110011110111;
		14'b10000010101000: color_data = 12'b110011110111;
		14'b10000010101001: color_data = 12'b110011110111;
		14'b10000010101010: color_data = 12'b110011110111;
		14'b10000010101011: color_data = 12'b110011110111;
		14'b10000010101100: color_data = 12'b110011110111;
		14'b10000010101101: color_data = 12'b110011110111;
		14'b10000010101110: color_data = 12'b110011110111;
		14'b10000010101111: color_data = 12'b110011110111;

		default: color_data = 12'b000000000000;
	endcase
endmodule
